-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity loader_firmware_rom is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end loader_firmware_rom;

architecture arch of loader_firmware_rom is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0ba9",
     9 => x"c4080b0b",
    10 => x"0ba9c808",
    11 => x"0b0b0ba9",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a9cc0c0b",
    16 => x"0b0ba9c8",
    17 => x"0c0b0b0b",
    18 => x"a9c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba0e8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a9c470ae",
    57 => x"f8278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"89d00402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"a9d40c9f",
    65 => x"0ba9d80c",
    66 => x"a0717081",
    67 => x"055334a9",
    68 => x"d808ff05",
    69 => x"a9d80ca9",
    70 => x"d8088025",
    71 => x"eb38a9d4",
    72 => x"08ff05a9",
    73 => x"d40ca9d4",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0ba9d4",
    94 => x"08258f38",
    95 => x"82b22da9",
    96 => x"d408ff05",
    97 => x"a9d40c82",
    98 => x"f404a9d4",
    99 => x"08a9d808",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38a9d408",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134a9",
   108 => x"d8088105",
   109 => x"a9d80ca9",
   110 => x"d808519f",
   111 => x"7125e238",
   112 => x"800ba9d8",
   113 => x"0ca9d408",
   114 => x"8105a9d4",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"a9d80881",
   120 => x"05a9d80c",
   121 => x"a9d808a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"a9d80ca9",
   125 => x"d4088105",
   126 => x"a9d40c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800ba9",
   155 => x"dc0cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820ba9dc",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"a9dc0884",
   167 => x"07a9dc0c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0ba6",
   172 => x"ac0c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2ca9dc08",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02d4050d",
   198 => x"a3e85185",
   199 => x"f32d97f8",
   200 => x"2da9c408",
   201 => x"802e81ef",
   202 => x"388ae72d",
   203 => x"a9c40853",
   204 => x"a9c40880",
   205 => x"2e81e238",
   206 => x"9abb2da9",
   207 => x"c408802e",
   208 => x"8738a480",
   209 => x"5186d504",
   210 => x"93e42da9",
   211 => x"c408802e",
   212 => x"8738a494",
   213 => x"5185f32d",
   214 => x"a4ac5185",
   215 => x"f32da4c0",
   216 => x"52a9e051",
   217 => x"90f92da9",
   218 => x"c408802e",
   219 => x"81a938a4",
   220 => x"cc5185f3",
   221 => x"2da9e408",
   222 => x"57807759",
   223 => x"5a767a2e",
   224 => x"8b38811a",
   225 => x"78812a59",
   226 => x"5a77f738",
   227 => x"f71a5a80",
   228 => x"772580fe",
   229 => x"38795277",
   230 => x"5184802d",
   231 => x"a9ec52a9",
   232 => x"e05193be",
   233 => x"2da9c408",
   234 => x"53a9c408",
   235 => x"802e80c9",
   236 => x"38a9ec5b",
   237 => x"805987e6",
   238 => x"047a7084",
   239 => x"055c0870",
   240 => x"81ff0671",
   241 => x"882c7081",
   242 => x"ff067390",
   243 => x"2c7081ff",
   244 => x"0675982a",
   245 => x"fec80cfe",
   246 => x"c80c58fe",
   247 => x"c80c57fe",
   248 => x"c80c841a",
   249 => x"5a537653",
   250 => x"84807725",
   251 => x"84388480",
   252 => x"53727924",
   253 => x"c4388882",
   254 => x"04a4dc51",
   255 => x"85f32d88",
   256 => x"9904a9e0",
   257 => x"5193912d",
   258 => x"fc801781",
   259 => x"19595787",
   260 => x"8f048153",
   261 => x"88990480",
   262 => x"5372a9c4",
   263 => x"0c02ac05",
   264 => x"0d0402f8",
   265 => x"050d9ef7",
   266 => x"2d81f72d",
   267 => x"815184e5",
   268 => x"2dfec452",
   269 => x"81720c9d",
   270 => x"c32d9dc3",
   271 => x"2d84720c",
   272 => x"73518694",
   273 => x"2da6f851",
   274 => x"a0d52d80",
   275 => x"5184e52d",
   276 => x"0288050d",
   277 => x"0402fc05",
   278 => x"0d825188",
   279 => x"a22d0284",
   280 => x"050d0402",
   281 => x"fc050d80",
   282 => x"5188a22d",
   283 => x"0284050d",
   284 => x"0402f405",
   285 => x"0d747081",
   286 => x"8432aee8",
   287 => x"0c708306",
   288 => x"525370a7",
   289 => x"d80b8805",
   290 => x"81b72d72",
   291 => x"892a7081",
   292 => x"06515170",
   293 => x"a8a80b81",
   294 => x"b72d7283",
   295 => x"2a810673",
   296 => x"882a7081",
   297 => x"06515252",
   298 => x"70802e85",
   299 => x"38718207",
   300 => x"5271a884",
   301 => x"0b81b72d",
   302 => x"72842c70",
   303 => x"83065151",
   304 => x"70a8900b",
   305 => x"81b72d70",
   306 => x"a9c40c02",
   307 => x"8c050d04",
   308 => x"02fc050d",
   309 => x"84b85188",
   310 => x"f12d810b",
   311 => x"fec40c84",
   312 => x"b80bfec0",
   313 => x"0c840bfe",
   314 => x"c40c830b",
   315 => x"fecc0c9d",
   316 => x"de2d9eeb",
   317 => x"2d9dc32d",
   318 => x"9dc32d81",
   319 => x"f72d8151",
   320 => x"84e52d9d",
   321 => x"c32d9dc3",
   322 => x"2d815184",
   323 => x"e52d8151",
   324 => x"86942da9",
   325 => x"c408802e",
   326 => x"8738a4ec",
   327 => x"518aa304",
   328 => x"a5805185",
   329 => x"f32d8a8e",
   330 => x"0402e805",
   331 => x"0d77797b",
   332 => x"58555580",
   333 => x"53727625",
   334 => x"a3387470",
   335 => x"81055680",
   336 => x"f52d7470",
   337 => x"81055680",
   338 => x"f52d5252",
   339 => x"71712e86",
   340 => x"3881518a",
   341 => x"de048113",
   342 => x"538ab504",
   343 => x"805170a9",
   344 => x"c40c0298",
   345 => x"050d0402",
   346 => x"d8050d80",
   347 => x"0badf40c",
   348 => x"a9ec5280",
   349 => x"5199a02d",
   350 => x"a9c40854",
   351 => x"a9c4088c",
   352 => x"38a59851",
   353 => x"85f32d73",
   354 => x"55908204",
   355 => x"8056810b",
   356 => x"ae980c88",
   357 => x"53a5a452",
   358 => x"aaa2518a",
   359 => x"a92da9c4",
   360 => x"08762e09",
   361 => x"81068738",
   362 => x"a9c408ae",
   363 => x"980c8853",
   364 => x"a5b052aa",
   365 => x"be518aa9",
   366 => x"2da9c408",
   367 => x"8738a9c4",
   368 => x"08ae980c",
   369 => x"ae980880",
   370 => x"2e80f638",
   371 => x"adb20b80",
   372 => x"f52dadb3",
   373 => x"0b80f52d",
   374 => x"71982b71",
   375 => x"902b07ad",
   376 => x"b40b80f5",
   377 => x"2d70882b",
   378 => x"7207adb5",
   379 => x"0b80f52d",
   380 => x"7107adea",
   381 => x"0b80f52d",
   382 => x"adeb0b80",
   383 => x"f52d7188",
   384 => x"2b07535f",
   385 => x"54525a56",
   386 => x"57557381",
   387 => x"abaa2e09",
   388 => x"81068d38",
   389 => x"75519ac2",
   390 => x"2da9c408",
   391 => x"568cad04",
   392 => x"7382d4d5",
   393 => x"2e8738a5",
   394 => x"bc518cee",
   395 => x"04a9ec52",
   396 => x"755199a0",
   397 => x"2da9c408",
   398 => x"55a9c408",
   399 => x"802e83c2",
   400 => x"388853a5",
   401 => x"b052aabe",
   402 => x"518aa92d",
   403 => x"a9c40889",
   404 => x"38810bad",
   405 => x"f40c8cf4",
   406 => x"048853a5",
   407 => x"a452aaa2",
   408 => x"518aa92d",
   409 => x"a9c40880",
   410 => x"2e8a38a5",
   411 => x"d05185f3",
   412 => x"2d8dce04",
   413 => x"adea0b80",
   414 => x"f52d5473",
   415 => x"80d52e09",
   416 => x"810680ca",
   417 => x"38adeb0b",
   418 => x"80f52d54",
   419 => x"7381aa2e",
   420 => x"098106ba",
   421 => x"38800ba9",
   422 => x"ec0b80f5",
   423 => x"2d565474",
   424 => x"81e92e83",
   425 => x"38815474",
   426 => x"81eb2e8c",
   427 => x"38805573",
   428 => x"752e0981",
   429 => x"0682cb38",
   430 => x"a9f70b80",
   431 => x"f52d5574",
   432 => x"8d38a9f8",
   433 => x"0b80f52d",
   434 => x"5473822e",
   435 => x"86388055",
   436 => x"908204a9",
   437 => x"f90b80f5",
   438 => x"2d70adec",
   439 => x"0cff05ad",
   440 => x"f00ca9fa",
   441 => x"0b80f52d",
   442 => x"a9fb0b80",
   443 => x"f52d5876",
   444 => x"05778280",
   445 => x"290570ad",
   446 => x"f80ca9fc",
   447 => x"0b80f52d",
   448 => x"70ae8c0c",
   449 => x"adf40859",
   450 => x"57587680",
   451 => x"2e81a338",
   452 => x"8853a5b0",
   453 => x"52aabe51",
   454 => x"8aa92da9",
   455 => x"c40881e2",
   456 => x"38adec08",
   457 => x"70842bae",
   458 => x"900c70ae",
   459 => x"880caa91",
   460 => x"0b80f52d",
   461 => x"aa900b80",
   462 => x"f52d7182",
   463 => x"802905aa",
   464 => x"920b80f5",
   465 => x"2d708480",
   466 => x"802912aa",
   467 => x"930b80f5",
   468 => x"2d708180",
   469 => x"0a291270",
   470 => x"ae940cae",
   471 => x"8c087129",
   472 => x"adf80805",
   473 => x"70adfc0c",
   474 => x"aa990b80",
   475 => x"f52daa98",
   476 => x"0b80f52d",
   477 => x"71828029",
   478 => x"05aa9a0b",
   479 => x"80f52d70",
   480 => x"84808029",
   481 => x"12aa9b0b",
   482 => x"80f52d70",
   483 => x"982b81f0",
   484 => x"0a067205",
   485 => x"70ae800c",
   486 => x"fe117e29",
   487 => x"7705ae84",
   488 => x"0c525952",
   489 => x"43545e51",
   490 => x"5259525d",
   491 => x"57595790",
   492 => x"8004a9fe",
   493 => x"0b80f52d",
   494 => x"a9fd0b80",
   495 => x"f52d7182",
   496 => x"80290570",
   497 => x"ae900c70",
   498 => x"a02983ff",
   499 => x"0570892a",
   500 => x"70ae880c",
   501 => x"aa830b80",
   502 => x"f52daa82",
   503 => x"0b80f52d",
   504 => x"71828029",
   505 => x"0570ae94",
   506 => x"0c7b7129",
   507 => x"1e70ae84",
   508 => x"0c7dae80",
   509 => x"0c7305ad",
   510 => x"fc0c555e",
   511 => x"51515555",
   512 => x"815574a9",
   513 => x"c40c02a8",
   514 => x"050d0402",
   515 => x"ec050d76",
   516 => x"70872c71",
   517 => x"80ff0655",
   518 => x"5654adf4",
   519 => x"088a3873",
   520 => x"882c7481",
   521 => x"ff065455",
   522 => x"a9ec52ad",
   523 => x"f8081551",
   524 => x"99a02da9",
   525 => x"c40854a9",
   526 => x"c408802e",
   527 => x"b338adf4",
   528 => x"08802e98",
   529 => x"38728429",
   530 => x"a9ec0570",
   531 => x"0852539a",
   532 => x"c22da9c4",
   533 => x"08f00a06",
   534 => x"5390ee04",
   535 => x"7210a9ec",
   536 => x"057080e0",
   537 => x"2d52539a",
   538 => x"f22da9c4",
   539 => x"08537254",
   540 => x"73a9c40c",
   541 => x"0294050d",
   542 => x"0402c805",
   543 => x"0d7f615f",
   544 => x"5b800bae",
   545 => x"8008ae84",
   546 => x"08595d56",
   547 => x"adf40876",
   548 => x"2e8a38ad",
   549 => x"ec08842b",
   550 => x"5891a204",
   551 => x"ae880884",
   552 => x"2b588059",
   553 => x"78782781",
   554 => x"a938788f",
   555 => x"06a01757",
   556 => x"54738f38",
   557 => x"a9ec5276",
   558 => x"51811757",
   559 => x"99a02da9",
   560 => x"ec568076",
   561 => x"80f52d56",
   562 => x"5474742e",
   563 => x"83388154",
   564 => x"7481e52e",
   565 => x"80f63881",
   566 => x"70750655",
   567 => x"5d73802e",
   568 => x"80ea388b",
   569 => x"1680f52d",
   570 => x"98065a79",
   571 => x"80de388b",
   572 => x"537d5275",
   573 => x"518aa92d",
   574 => x"a9c40880",
   575 => x"cf389c16",
   576 => x"08519ac2",
   577 => x"2da9c408",
   578 => x"841c0c9a",
   579 => x"1680e02d",
   580 => x"519af22d",
   581 => x"a9c408a9",
   582 => x"c408881d",
   583 => x"0ca9c408",
   584 => x"5555adf4",
   585 => x"08802e98",
   586 => x"38941680",
   587 => x"e02d519a",
   588 => x"f22da9c4",
   589 => x"08902b83",
   590 => x"fff00a06",
   591 => x"70165154",
   592 => x"73881c0c",
   593 => x"797b0c7c",
   594 => x"54938804",
   595 => x"81195991",
   596 => x"a404adf4",
   597 => x"08802eae",
   598 => x"387b5190",
   599 => x"8b2da9c4",
   600 => x"08a9c408",
   601 => x"80ffffff",
   602 => x"f806555c",
   603 => x"7380ffff",
   604 => x"fff82e92",
   605 => x"38a9c408",
   606 => x"fe05adec",
   607 => x"0829adfc",
   608 => x"08055791",
   609 => x"a2048054",
   610 => x"73a9c40c",
   611 => x"02b8050d",
   612 => x"0402f405",
   613 => x"0d747008",
   614 => x"8105710c",
   615 => x"7008adf0",
   616 => x"08065353",
   617 => x"718e3888",
   618 => x"13085190",
   619 => x"8b2da9c4",
   620 => x"0888140c",
   621 => x"810ba9c4",
   622 => x"0c028c05",
   623 => x"0d0402f0",
   624 => x"050d7588",
   625 => x"1108fe05",
   626 => x"adec0829",
   627 => x"adfc0811",
   628 => x"7208adf0",
   629 => x"08060579",
   630 => x"55535454",
   631 => x"99a02d02",
   632 => x"90050d04",
   633 => x"adf408a9",
   634 => x"c40c0402",
   635 => x"f4050dd4",
   636 => x"5281ff72",
   637 => x"0c710853",
   638 => x"81ff720c",
   639 => x"72882b83",
   640 => x"fe800672",
   641 => x"087081ff",
   642 => x"06515253",
   643 => x"81ff720c",
   644 => x"72710788",
   645 => x"2b720870",
   646 => x"81ff0651",
   647 => x"525381ff",
   648 => x"720c7271",
   649 => x"07882b72",
   650 => x"087081ff",
   651 => x"067207a9",
   652 => x"c40c5253",
   653 => x"028c050d",
   654 => x"0402f405",
   655 => x"0d747671",
   656 => x"81ff06d4",
   657 => x"0c5353ae",
   658 => x"9c088538",
   659 => x"71892b52",
   660 => x"71982ad4",
   661 => x"0c71902a",
   662 => x"7081ff06",
   663 => x"d40c5171",
   664 => x"882a7081",
   665 => x"ff06d40c",
   666 => x"517181ff",
   667 => x"06d40c72",
   668 => x"902a7081",
   669 => x"ff06d40c",
   670 => x"51d40870",
   671 => x"81ff0651",
   672 => x"5182b8bf",
   673 => x"527081ff",
   674 => x"2e098106",
   675 => x"943881ff",
   676 => x"0bd40cd4",
   677 => x"087081ff",
   678 => x"06ff1454",
   679 => x"515171e5",
   680 => x"3870a9c4",
   681 => x"0c028c05",
   682 => x"0d0402fc",
   683 => x"050d81c7",
   684 => x"5181ff0b",
   685 => x"d40cff11",
   686 => x"51708025",
   687 => x"f4380284",
   688 => x"050d0402",
   689 => x"f0050d95",
   690 => x"aa2d8fcf",
   691 => x"53805287",
   692 => x"fc80f751",
   693 => x"94b92da9",
   694 => x"c40854a9",
   695 => x"c408812e",
   696 => x"098106a3",
   697 => x"3881ff0b",
   698 => x"d40c820a",
   699 => x"52849c80",
   700 => x"e95194b9",
   701 => x"2da9c408",
   702 => x"8b3881ff",
   703 => x"0bd40c73",
   704 => x"53968d04",
   705 => x"95aa2dff",
   706 => x"135372c1",
   707 => x"3872a9c4",
   708 => x"0c029005",
   709 => x"0d0402f4",
   710 => x"050d81ff",
   711 => x"0bd40c93",
   712 => x"53805287",
   713 => x"fc80c151",
   714 => x"94b92da9",
   715 => x"c4088b38",
   716 => x"81ff0bd4",
   717 => x"0c815396",
   718 => x"c30495aa",
   719 => x"2dff1353",
   720 => x"72df3872",
   721 => x"a9c40c02",
   722 => x"8c050d04",
   723 => x"02f0050d",
   724 => x"95aa2d83",
   725 => x"aa52849c",
   726 => x"80c85194",
   727 => x"b92da9c4",
   728 => x"08812e09",
   729 => x"81069238",
   730 => x"93eb2da9",
   731 => x"c40883ff",
   732 => x"ff065372",
   733 => x"83aa2e97",
   734 => x"3896962d",
   735 => x"978a0481",
   736 => x"5497ef04",
   737 => x"a5dc5185",
   738 => x"f32d8054",
   739 => x"97ef0481",
   740 => x"ff0bd40c",
   741 => x"b15395c3",
   742 => x"2da9c408",
   743 => x"802e80c0",
   744 => x"38805287",
   745 => x"fc80fa51",
   746 => x"94b92da9",
   747 => x"c408b138",
   748 => x"81ff0bd4",
   749 => x"0cd40853",
   750 => x"81ff0bd4",
   751 => x"0c81ff0b",
   752 => x"d40c81ff",
   753 => x"0bd40c81",
   754 => x"ff0bd40c",
   755 => x"72862a70",
   756 => x"8106a9c4",
   757 => x"08565153",
   758 => x"72802e93",
   759 => x"3896ff04",
   760 => x"72822eff",
   761 => x"9f38ff13",
   762 => x"5372ffaa",
   763 => x"38725473",
   764 => x"a9c40c02",
   765 => x"90050d04",
   766 => x"02f0050d",
   767 => x"810bae9c",
   768 => x"0c8454d0",
   769 => x"08708f2a",
   770 => x"70810651",
   771 => x"515372f3",
   772 => x"3872d00c",
   773 => x"95aa2da5",
   774 => x"ec5185f3",
   775 => x"2dd00870",
   776 => x"8f2a7081",
   777 => x"06515153",
   778 => x"72f33881",
   779 => x"0bd00cb1",
   780 => x"53805284",
   781 => x"d480c051",
   782 => x"94b92da9",
   783 => x"c408812e",
   784 => x"a1387282",
   785 => x"2e098106",
   786 => x"8c38a5f8",
   787 => x"5185f32d",
   788 => x"80539997",
   789 => x"04ff1353",
   790 => x"72d738ff",
   791 => x"145473ff",
   792 => x"a23896cc",
   793 => x"2da9c408",
   794 => x"ae9c0ca9",
   795 => x"c4088b38",
   796 => x"815287fc",
   797 => x"80d05194",
   798 => x"b92d81ff",
   799 => x"0bd40cd0",
   800 => x"08708f2a",
   801 => x"70810651",
   802 => x"515372f3",
   803 => x"3872d00c",
   804 => x"81ff0bd4",
   805 => x"0c815372",
   806 => x"a9c40c02",
   807 => x"90050d04",
   808 => x"02e8050d",
   809 => x"78558056",
   810 => x"81ff0bd4",
   811 => x"0cd00870",
   812 => x"8f2a7081",
   813 => x"06515153",
   814 => x"72f33882",
   815 => x"810bd00c",
   816 => x"81ff0bd4",
   817 => x"0c775287",
   818 => x"fc80d151",
   819 => x"94b92d80",
   820 => x"dbc6df54",
   821 => x"a9c40880",
   822 => x"2e8a38a4",
   823 => x"dc5185f3",
   824 => x"2d9ab204",
   825 => x"81ff0bd4",
   826 => x"0cd40870",
   827 => x"81ff0651",
   828 => x"537281fe",
   829 => x"2e098106",
   830 => x"9d3880ff",
   831 => x"5393eb2d",
   832 => x"a9c40875",
   833 => x"70840557",
   834 => x"0cff1353",
   835 => x"728025ed",
   836 => x"3881569a",
   837 => x"9c04ff14",
   838 => x"5473c938",
   839 => x"81ff0bd4",
   840 => x"0cd00870",
   841 => x"8f2a7081",
   842 => x"06515153",
   843 => x"72f33872",
   844 => x"d00c75a9",
   845 => x"c40c0298",
   846 => x"050d04ae",
   847 => x"9c08a9c4",
   848 => x"0c0402f4",
   849 => x"050d7470",
   850 => x"882a83fe",
   851 => x"80067072",
   852 => x"982a0772",
   853 => x"882b87fc",
   854 => x"80800673",
   855 => x"982b81f0",
   856 => x"0a067173",
   857 => x"0707a9c4",
   858 => x"0c565153",
   859 => x"51028c05",
   860 => x"0d0402f8",
   861 => x"050d028e",
   862 => x"0580f52d",
   863 => x"74882b07",
   864 => x"7083ffff",
   865 => x"06a9c40c",
   866 => x"51028805",
   867 => x"0d0402fc",
   868 => x"050d7251",
   869 => x"80710c80",
   870 => x"0b84120c",
   871 => x"0284050d",
   872 => x"0402f405",
   873 => x"0d9ef12d",
   874 => x"e008e408",
   875 => x"718b2a70",
   876 => x"81065153",
   877 => x"54527080",
   878 => x"2e9d38ae",
   879 => x"a0087084",
   880 => x"29aea805",
   881 => x"7381ff06",
   882 => x"710c5151",
   883 => x"aea00881",
   884 => x"118706ae",
   885 => x"a00c5172",
   886 => x"8b2a7081",
   887 => x"06515170",
   888 => x"802e8192",
   889 => x"38a8fc08",
   890 => x"8429aed4",
   891 => x"057381ff",
   892 => x"06710c51",
   893 => x"a8fc0881",
   894 => x"05a8fc0c",
   895 => x"850ba8f8",
   896 => x"0ca8fc08",
   897 => x"a8f4082e",
   898 => x"09810681",
   899 => x"a638800b",
   900 => x"a8fc0cae",
   901 => x"e408819b",
   902 => x"38aed408",
   903 => x"70097083",
   904 => x"06fecc0c",
   905 => x"5270852a",
   906 => x"708106ae",
   907 => x"cc085551",
   908 => x"52537080",
   909 => x"2e8e38ae",
   910 => x"dc08fe80",
   911 => x"3212aecc",
   912 => x"0c9ccb04",
   913 => x"aedc0812",
   914 => x"aecc0c72",
   915 => x"842a7081",
   916 => x"06aec808",
   917 => x"54515170",
   918 => x"802e9038",
   919 => x"aed80881",
   920 => x"ff321281",
   921 => x"05aec80c",
   922 => x"9db30471",
   923 => x"aed80831",
   924 => x"aec80c9d",
   925 => x"b304a8f8",
   926 => x"08ff05a8",
   927 => x"f80ca8f8",
   928 => x"08ff2e09",
   929 => x"8106ac38",
   930 => x"a8fc0880",
   931 => x"2e923881",
   932 => x"0baee40c",
   933 => x"870ba8f4",
   934 => x"0831a8f4",
   935 => x"0c9dae04",
   936 => x"aee40851",
   937 => x"70802e86",
   938 => x"38ff11ae",
   939 => x"e40c800b",
   940 => x"a8fc0c80",
   941 => x"0baed00c",
   942 => x"9ee42d9e",
   943 => x"eb2d028c",
   944 => x"050d0402",
   945 => x"fc050d9e",
   946 => x"f12d810b",
   947 => x"aed00c9e",
   948 => x"eb2daed0",
   949 => x"085170fa",
   950 => x"38028405",
   951 => x"0d0402f8",
   952 => x"050daea0",
   953 => x"519b8e2d",
   954 => x"800baee4",
   955 => x"0c830ba8",
   956 => x"f40ce408",
   957 => x"708c2a70",
   958 => x"81065151",
   959 => x"5271802e",
   960 => x"8638840b",
   961 => x"a8f40ce4",
   962 => x"08708d2a",
   963 => x"70810651",
   964 => x"51527180",
   965 => x"2e9f3887",
   966 => x"0ba8f408",
   967 => x"31a8f40c",
   968 => x"e408708a",
   969 => x"2a708106",
   970 => x"51515271",
   971 => x"802ef138",
   972 => x"81f40be4",
   973 => x"0c9ba151",
   974 => x"9ee02d9e",
   975 => x"c32d0288",
   976 => x"050d0402",
   977 => x"f8050da9",
   978 => x"80528f51",
   979 => x"80727084",
   980 => x"05540cff",
   981 => x"11517080",
   982 => x"25f23802",
   983 => x"88050d04",
   984 => x"71980c04",
   985 => x"ffb008a9",
   986 => x"c40c0481",
   987 => x"0bffb00c",
   988 => x"04800bff",
   989 => x"b00c0402",
   990 => x"fc050d80",
   991 => x"0ba9c00c",
   992 => x"805184e5",
   993 => x"2d028405",
   994 => x"0d0402ec",
   995 => x"050d7654",
   996 => x"8052870b",
   997 => x"881580f5",
   998 => x"2d565374",
   999 => x"72248338",
  1000 => x"a0537251",
  1001 => x"82ee2d81",
  1002 => x"128b1580",
  1003 => x"f52d5452",
  1004 => x"727225de",
  1005 => x"38029405",
  1006 => x"0d0402f0",
  1007 => x"050daeec",
  1008 => x"085481f7",
  1009 => x"2d800bae",
  1010 => x"f00c7308",
  1011 => x"802e8180",
  1012 => x"38820ba9",
  1013 => x"d80caef0",
  1014 => x"088f06a9",
  1015 => x"d40c7308",
  1016 => x"5271832e",
  1017 => x"96387183",
  1018 => x"26893871",
  1019 => x"812eaf38",
  1020 => x"a0bb0471",
  1021 => x"852e9f38",
  1022 => x"a0bb0488",
  1023 => x"1480f52d",
  1024 => x"841508a6",
  1025 => x"a0535452",
  1026 => x"85f32d71",
  1027 => x"84291370",
  1028 => x"085252a0",
  1029 => x"bf047351",
  1030 => x"9f8a2da0",
  1031 => x"bb04aee8",
  1032 => x"08881508",
  1033 => x"2c708106",
  1034 => x"51527180",
  1035 => x"2e8738a6",
  1036 => x"a451a0b8",
  1037 => x"04a6a851",
  1038 => x"85f32d84",
  1039 => x"14085185",
  1040 => x"f32daef0",
  1041 => x"088105ae",
  1042 => x"f00c8c14",
  1043 => x"549fca04",
  1044 => x"0290050d",
  1045 => x"0471aeec",
  1046 => x"0c9fba2d",
  1047 => x"aef008ff",
  1048 => x"05aef40c",
  1049 => x"04000000",
  1050 => x"00ffffff",
  1051 => x"ff00ffff",
  1052 => x"ffff00ff",
  1053 => x"ffffff00",
  1054 => x"4d617374",
  1055 => x"65720000",
  1056 => x"4f504c4c",
  1057 => x"00000000",
  1058 => x"53434300",
  1059 => x"50534700",
  1060 => x"4261636b",
  1061 => x"00000000",
  1062 => x"52657365",
  1063 => x"74000000",
  1064 => x"53617665",
  1065 => x"20616e64",
  1066 => x"20526573",
  1067 => x"65740000",
  1068 => x"4f707469",
  1069 => x"6f6e7320",
  1070 => x"10000000",
  1071 => x"536f756e",
  1072 => x"64201000",
  1073 => x"54757262",
  1074 => x"6f000000",
  1075 => x"4d6f7573",
  1076 => x"6520656d",
  1077 => x"756c6174",
  1078 => x"696f6e00",
  1079 => x"45786974",
  1080 => x"00000000",
  1081 => x"5363616e",
  1082 => x"6c696e65",
  1083 => x"73000000",
  1084 => x"53442043",
  1085 => x"61726400",
  1086 => x"4a617061",
  1087 => x"6e657365",
  1088 => x"206b6579",
  1089 => x"206c6179",
  1090 => x"6f757400",
  1091 => x"32303438",
  1092 => x"4b422052",
  1093 => x"414d0000",
  1094 => x"34303936",
  1095 => x"4b422052",
  1096 => x"414d0000",
  1097 => x"536c323a",
  1098 => x"204e6f6e",
  1099 => x"65000000",
  1100 => x"536c323a",
  1101 => x"20455345",
  1102 => x"2d534343",
  1103 => x"20314d42",
  1104 => x"2f534343",
  1105 => x"2d490000",
  1106 => x"536c323a",
  1107 => x"20455345",
  1108 => x"2d52414d",
  1109 => x"20314d42",
  1110 => x"2f415343",
  1111 => x"49493800",
  1112 => x"536c323a",
  1113 => x"20455345",
  1114 => x"2d52414d",
  1115 => x"20314d42",
  1116 => x"2f415343",
  1117 => x"49493136",
  1118 => x"00000000",
  1119 => x"536c313a",
  1120 => x"204e6f6e",
  1121 => x"65000000",
  1122 => x"536c313a",
  1123 => x"20455345",
  1124 => x"2d534343",
  1125 => x"20314d42",
  1126 => x"2f534343",
  1127 => x"2d490000",
  1128 => x"536c313a",
  1129 => x"204d6567",
  1130 => x"6152414d",
  1131 => x"00000000",
  1132 => x"56474120",
  1133 => x"2d203331",
  1134 => x"4b487a2c",
  1135 => x"20363048",
  1136 => x"7a000000",
  1137 => x"56474120",
  1138 => x"2d203331",
  1139 => x"4b487a2c",
  1140 => x"20353048",
  1141 => x"7a000000",
  1142 => x"5456202d",
  1143 => x"20343830",
  1144 => x"692c2036",
  1145 => x"30487a00",
  1146 => x"496e6974",
  1147 => x"69616c69",
  1148 => x"7a696e67",
  1149 => x"20534420",
  1150 => x"63617264",
  1151 => x"0a000000",
  1152 => x"53444843",
  1153 => x"20636172",
  1154 => x"64206465",
  1155 => x"74656374",
  1156 => x"65640a00",
  1157 => x"46617433",
  1158 => x"32206e6f",
  1159 => x"74207375",
  1160 => x"70706f72",
  1161 => x"7465640a",
  1162 => x"00000000",
  1163 => x"54727969",
  1164 => x"6e672053",
  1165 => x"50454343",
  1166 => x"592e524f",
  1167 => x"4d0a0000",
  1168 => x"53504543",
  1169 => x"43592020",
  1170 => x"524f4d00",
  1171 => x"4c6f6164",
  1172 => x"696e6720",
  1173 => x"42494f53",
  1174 => x"0a000000",
  1175 => x"52656164",
  1176 => x"20666169",
  1177 => x"6c65640a",
  1178 => x"00000000",
  1179 => x"4c6f6164",
  1180 => x"696e6720",
  1181 => x"42494f53",
  1182 => x"20646f6e",
  1183 => x"650a0000",
  1184 => x"4c6f6164",
  1185 => x"696e6720",
  1186 => x"42494f53",
  1187 => x"20666169",
  1188 => x"6c65640a",
  1189 => x"00000000",
  1190 => x"4d425220",
  1191 => x"6661696c",
  1192 => x"0a000000",
  1193 => x"46415431",
  1194 => x"36202020",
  1195 => x"00000000",
  1196 => x"46415433",
  1197 => x"32202020",
  1198 => x"00000000",
  1199 => x"4e6f2070",
  1200 => x"61727469",
  1201 => x"74696f6e",
  1202 => x"20736967",
  1203 => x"0a000000",
  1204 => x"42616420",
  1205 => x"70617274",
  1206 => x"0a000000",
  1207 => x"53444843",
  1208 => x"20657272",
  1209 => x"6f72210a",
  1210 => x"00000000",
  1211 => x"53442069",
  1212 => x"6e69742e",
  1213 => x"2e2e0a00",
  1214 => x"53442063",
  1215 => x"61726420",
  1216 => x"72657365",
  1217 => x"74206661",
  1218 => x"696c6564",
  1219 => x"210a0000",
  1220 => x"57726974",
  1221 => x"65206661",
  1222 => x"696c6564",
  1223 => x"0a000000",
  1224 => x"16200000",
  1225 => x"14200000",
  1226 => x"15200000",
  1227 => x"00000002",
  1228 => x"00000005",
  1229 => x"00001078",
  1230 => x"00000007",
  1231 => x"00000005",
  1232 => x"00001080",
  1233 => x"00000007",
  1234 => x"00000005",
  1235 => x"00001088",
  1236 => x"00000007",
  1237 => x"00000005",
  1238 => x"0000108c",
  1239 => x"00000007",
  1240 => x"00000004",
  1241 => x"00001090",
  1242 => x"00001378",
  1243 => x"00000000",
  1244 => x"00000000",
  1245 => x"00000000",
  1246 => x"00000002",
  1247 => x"00001098",
  1248 => x"00000463",
  1249 => x"00000002",
  1250 => x"000010a0",
  1251 => x"00000455",
  1252 => x"00000004",
  1253 => x"000010b0",
  1254 => x"000013d8",
  1255 => x"00000004",
  1256 => x"000010bc",
  1257 => x"00001330",
  1258 => x"00000001",
  1259 => x"000010c4",
  1260 => x"00000007",
  1261 => x"00000001",
  1262 => x"000010cc",
  1263 => x"0000000a",
  1264 => x"00000002",
  1265 => x"000010dc",
  1266 => x"00000f77",
  1267 => x"00000000",
  1268 => x"00000000",
  1269 => x"00000000",
  1270 => x"00000003",
  1271 => x"00001468",
  1272 => x"00000003",
  1273 => x"00000001",
  1274 => x"000010e4",
  1275 => x"0000000b",
  1276 => x"00000001",
  1277 => x"000010f0",
  1278 => x"00000002",
  1279 => x"00000003",
  1280 => x"0000145c",
  1281 => x"00000003",
  1282 => x"00000003",
  1283 => x"0000144c",
  1284 => x"00000004",
  1285 => x"00000001",
  1286 => x"000010f8",
  1287 => x"00000006",
  1288 => x"00000003",
  1289 => x"00001444",
  1290 => x"00000002",
  1291 => x"00000004",
  1292 => x"00001090",
  1293 => x"00001378",
  1294 => x"00000000",
  1295 => x"00000000",
  1296 => x"00000000",
  1297 => x"0000110c",
  1298 => x"00001118",
  1299 => x"00001124",
  1300 => x"00001130",
  1301 => x"00001148",
  1302 => x"00001160",
  1303 => x"0000117c",
  1304 => x"00001188",
  1305 => x"000011a0",
  1306 => x"000011b0",
  1307 => x"000011c4",
  1308 => x"000011d8",
  1309 => x"00000003",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

