-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity loader_firmware_rom is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end loader_firmware_rom;

architecture arch of loader_firmware_rom is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0ba0",
     9 => x"c0080b0b",
    10 => x"0ba0c408",
    11 => x"0b0b0ba0",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a0c80c0b",
    16 => x"0b0ba0c4",
    17 => x"0c0b0b0b",
    18 => x"a0c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0b9dac",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a0c070a5",
    57 => x"e4278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"86940402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"a0d00c9f",
    65 => x"0ba0d40c",
    66 => x"a0717081",
    67 => x"055334a0",
    68 => x"d408ff05",
    69 => x"a0d40ca0",
    70 => x"d4088025",
    71 => x"eb38a0d0",
    72 => x"08ff05a0",
    73 => x"d00ca0d0",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0ba0d0",
    94 => x"08258f38",
    95 => x"82b22da0",
    96 => x"d008ff05",
    97 => x"a0d00c82",
    98 => x"f404a0d0",
    99 => x"08a0d408",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38a0d008",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134a0",
   108 => x"d4088105",
   109 => x"a0d40ca0",
   110 => x"d408519f",
   111 => x"7125e238",
   112 => x"800ba0d4",
   113 => x"0ca0d008",
   114 => x"8105a0d0",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"a0d40881",
   120 => x"05a0d40c",
   121 => x"a0d408a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"a0d40ca0",
   125 => x"d0088105",
   126 => x"a0d00c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800ba0",
   155 => x"d80cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820ba0d8",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"a0d80884",
   167 => x"07a0d80c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0b9f",
   172 => x"f00c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2ca0d808",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02d4050d",
   198 => x"810bfec4",
   199 => x"0c840bfe",
   200 => x"c40c830b",
   201 => x"fecc0c9c",
   202 => x"902d9d9d",
   203 => x"2d9bf52d",
   204 => x"9bf52d81",
   205 => x"f72d8151",
   206 => x"84e52d9b",
   207 => x"f52d9bf5",
   208 => x"2d80ff53",
   209 => x"9bf52d81",
   210 => x"5184e52d",
   211 => x"ff135372",
   212 => x"8025f138",
   213 => x"9bf52d9b",
   214 => x"f52d9dbc",
   215 => x"5185f32d",
   216 => x"96aa2da0",
   217 => x"c008802e",
   218 => x"81e83889",
   219 => x"992da0c0",
   220 => x"08802e81",
   221 => x"dd3898ed",
   222 => x"2da0c008",
   223 => x"802e8738",
   224 => x"9dd45185",
   225 => x"f32d9296",
   226 => x"2da0c008",
   227 => x"802e8738",
   228 => x"9de85185",
   229 => x"f32d9df8",
   230 => x"5185f32d",
   231 => x"9e8c52a0",
   232 => x"dc518fab",
   233 => x"2da0c008",
   234 => x"802e81a6",
   235 => x"389e9851",
   236 => x"85f32da0",
   237 => x"e0085780",
   238 => x"77595a76",
   239 => x"7a2e8b38",
   240 => x"811a7881",
   241 => x"2a595a77",
   242 => x"f738f71a",
   243 => x"5a807725",
   244 => x"80fa3879",
   245 => x"52775184",
   246 => x"802da0e8",
   247 => x"52a0dc51",
   248 => x"91f02da0",
   249 => x"c008802e",
   250 => x"80c938a0",
   251 => x"e85b8059",
   252 => x"88a0047a",
   253 => x"7084055c",
   254 => x"087081ff",
   255 => x"0671882c",
   256 => x"7081ff06",
   257 => x"73902c70",
   258 => x"81ff0675",
   259 => x"982afec8",
   260 => x"0cfec80c",
   261 => x"58fec80c",
   262 => x"57fec80c",
   263 => x"841a5a53",
   264 => x"76538480",
   265 => x"77258438",
   266 => x"84805372",
   267 => x"7924c438",
   268 => x"88bc049e",
   269 => x"ac5185f3",
   270 => x"2d88d204",
   271 => x"a0dc5191",
   272 => x"c32dfc80",
   273 => x"17811959",
   274 => x"5787cd04",
   275 => x"9ebc5188",
   276 => x"d5049ed0",
   277 => x"5185f32d",
   278 => x"86da0402",
   279 => x"e8050d77",
   280 => x"797b5855",
   281 => x"55805372",
   282 => x"7625a338",
   283 => x"74708105",
   284 => x"5680f52d",
   285 => x"74708105",
   286 => x"5680f52d",
   287 => x"52527171",
   288 => x"2e863881",
   289 => x"51899004",
   290 => x"81135388",
   291 => x"e7048051",
   292 => x"70a0c00c",
   293 => x"0298050d",
   294 => x"0402d805",
   295 => x"0d800ba4",
   296 => x"f00ca0e8",
   297 => x"52805197",
   298 => x"d22da0c0",
   299 => x"0854a0c0",
   300 => x"088c389e",
   301 => x"e85185f3",
   302 => x"2d73558e",
   303 => x"b4048056",
   304 => x"810ba594",
   305 => x"0c88539e",
   306 => x"f452a19e",
   307 => x"5188db2d",
   308 => x"a0c00876",
   309 => x"2e098106",
   310 => x"8738a0c0",
   311 => x"08a5940c",
   312 => x"88539f80",
   313 => x"52a1ba51",
   314 => x"88db2da0",
   315 => x"c0088738",
   316 => x"a0c008a5",
   317 => x"940ca594",
   318 => x"08802e80",
   319 => x"f638a4ae",
   320 => x"0b80f52d",
   321 => x"a4af0b80",
   322 => x"f52d7198",
   323 => x"2b71902b",
   324 => x"07a4b00b",
   325 => x"80f52d70",
   326 => x"882b7207",
   327 => x"a4b10b80",
   328 => x"f52d7107",
   329 => x"a4e60b80",
   330 => x"f52da4e7",
   331 => x"0b80f52d",
   332 => x"71882b07",
   333 => x"535f5452",
   334 => x"5a565755",
   335 => x"7381abaa",
   336 => x"2e098106",
   337 => x"8d387551",
   338 => x"98f42da0",
   339 => x"c008568a",
   340 => x"df047382",
   341 => x"d4d52e87",
   342 => x"389f8c51",
   343 => x"8ba004a0",
   344 => x"e8527551",
   345 => x"97d22da0",
   346 => x"c00855a0",
   347 => x"c008802e",
   348 => x"83c23888",
   349 => x"539f8052",
   350 => x"a1ba5188",
   351 => x"db2da0c0",
   352 => x"08893881",
   353 => x"0ba4f00c",
   354 => x"8ba60488",
   355 => x"539ef452",
   356 => x"a19e5188",
   357 => x"db2da0c0",
   358 => x"08802e8a",
   359 => x"389fa051",
   360 => x"85f32d8c",
   361 => x"8004a4e6",
   362 => x"0b80f52d",
   363 => x"547380d5",
   364 => x"2e098106",
   365 => x"80ca38a4",
   366 => x"e70b80f5",
   367 => x"2d547381",
   368 => x"aa2e0981",
   369 => x"06ba3880",
   370 => x"0ba0e80b",
   371 => x"80f52d56",
   372 => x"547481e9",
   373 => x"2e833881",
   374 => x"547481eb",
   375 => x"2e8c3880",
   376 => x"5573752e",
   377 => x"09810682",
   378 => x"cb38a0f3",
   379 => x"0b80f52d",
   380 => x"55748d38",
   381 => x"a0f40b80",
   382 => x"f52d5473",
   383 => x"822e8638",
   384 => x"80558eb4",
   385 => x"04a0f50b",
   386 => x"80f52d70",
   387 => x"a4e80cff",
   388 => x"05a4ec0c",
   389 => x"a0f60b80",
   390 => x"f52da0f7",
   391 => x"0b80f52d",
   392 => x"58760577",
   393 => x"82802905",
   394 => x"70a4f40c",
   395 => x"a0f80b80",
   396 => x"f52d70a5",
   397 => x"880ca4f0",
   398 => x"08595758",
   399 => x"76802e81",
   400 => x"a3388853",
   401 => x"9f8052a1",
   402 => x"ba5188db",
   403 => x"2da0c008",
   404 => x"81e238a4",
   405 => x"e8087084",
   406 => x"2ba58c0c",
   407 => x"70a5840c",
   408 => x"a18d0b80",
   409 => x"f52da18c",
   410 => x"0b80f52d",
   411 => x"71828029",
   412 => x"05a18e0b",
   413 => x"80f52d70",
   414 => x"84808029",
   415 => x"12a18f0b",
   416 => x"80f52d70",
   417 => x"81800a29",
   418 => x"1270a590",
   419 => x"0ca58808",
   420 => x"7129a4f4",
   421 => x"080570a4",
   422 => x"f80ca195",
   423 => x"0b80f52d",
   424 => x"a1940b80",
   425 => x"f52d7182",
   426 => x"802905a1",
   427 => x"960b80f5",
   428 => x"2d708480",
   429 => x"802912a1",
   430 => x"970b80f5",
   431 => x"2d70982b",
   432 => x"81f00a06",
   433 => x"720570a4",
   434 => x"fc0cfe11",
   435 => x"7e297705",
   436 => x"a5800c52",
   437 => x"59524354",
   438 => x"5e515259",
   439 => x"525d5759",
   440 => x"578eb204",
   441 => x"a0fa0b80",
   442 => x"f52da0f9",
   443 => x"0b80f52d",
   444 => x"71828029",
   445 => x"0570a58c",
   446 => x"0c70a029",
   447 => x"83ff0570",
   448 => x"892a70a5",
   449 => x"840ca0ff",
   450 => x"0b80f52d",
   451 => x"a0fe0b80",
   452 => x"f52d7182",
   453 => x"80290570",
   454 => x"a5900c7b",
   455 => x"71291e70",
   456 => x"a5800c7d",
   457 => x"a4fc0c73",
   458 => x"05a4f80c",
   459 => x"555e5151",
   460 => x"55558155",
   461 => x"74a0c00c",
   462 => x"02a8050d",
   463 => x"0402ec05",
   464 => x"0d767087",
   465 => x"2c7180ff",
   466 => x"06555654",
   467 => x"a4f0088a",
   468 => x"3873882c",
   469 => x"7481ff06",
   470 => x"5455a0e8",
   471 => x"52a4f408",
   472 => x"155197d2",
   473 => x"2da0c008",
   474 => x"54a0c008",
   475 => x"802eb338",
   476 => x"a4f00880",
   477 => x"2e983872",
   478 => x"8429a0e8",
   479 => x"05700852",
   480 => x"5398f42d",
   481 => x"a0c008f0",
   482 => x"0a06538f",
   483 => x"a0047210",
   484 => x"a0e80570",
   485 => x"80e02d52",
   486 => x"5399a42d",
   487 => x"a0c00853",
   488 => x"725473a0",
   489 => x"c00c0294",
   490 => x"050d0402",
   491 => x"c8050d7f",
   492 => x"615f5b80",
   493 => x"0ba4fc08",
   494 => x"a5800859",
   495 => x"5d56a4f0",
   496 => x"08762e8a",
   497 => x"38a4e808",
   498 => x"842b588f",
   499 => x"d404a584",
   500 => x"08842b58",
   501 => x"80597878",
   502 => x"2781a938",
   503 => x"788f06a0",
   504 => x"17575473",
   505 => x"8f38a0e8",
   506 => x"52765181",
   507 => x"175797d2",
   508 => x"2da0e856",
   509 => x"807680f5",
   510 => x"2d565474",
   511 => x"742e8338",
   512 => x"81547481",
   513 => x"e52e80f6",
   514 => x"38817075",
   515 => x"06555d73",
   516 => x"802e80ea",
   517 => x"388b1680",
   518 => x"f52d9806",
   519 => x"5a7980de",
   520 => x"388b537d",
   521 => x"52755188",
   522 => x"db2da0c0",
   523 => x"0880cf38",
   524 => x"9c160851",
   525 => x"98f42da0",
   526 => x"c008841c",
   527 => x"0c9a1680",
   528 => x"e02d5199",
   529 => x"a42da0c0",
   530 => x"08a0c008",
   531 => x"881d0ca0",
   532 => x"c0085555",
   533 => x"a4f00880",
   534 => x"2e983894",
   535 => x"1680e02d",
   536 => x"5199a42d",
   537 => x"a0c00890",
   538 => x"2b83fff0",
   539 => x"0a067016",
   540 => x"51547388",
   541 => x"1c0c797b",
   542 => x"0c7c5491",
   543 => x"ba048119",
   544 => x"598fd604",
   545 => x"a4f00880",
   546 => x"2eae387b",
   547 => x"518ebd2d",
   548 => x"a0c008a0",
   549 => x"c00880ff",
   550 => x"fffff806",
   551 => x"555c7380",
   552 => x"fffffff8",
   553 => x"2e9238a0",
   554 => x"c008fe05",
   555 => x"a4e80829",
   556 => x"a4f80805",
   557 => x"578fd404",
   558 => x"805473a0",
   559 => x"c00c02b8",
   560 => x"050d0402",
   561 => x"f4050d74",
   562 => x"70088105",
   563 => x"710c7008",
   564 => x"a4ec0806",
   565 => x"5353718e",
   566 => x"38881308",
   567 => x"518ebd2d",
   568 => x"a0c00888",
   569 => x"140c810b",
   570 => x"a0c00c02",
   571 => x"8c050d04",
   572 => x"02f0050d",
   573 => x"75881108",
   574 => x"fe05a4e8",
   575 => x"0829a4f8",
   576 => x"08117208",
   577 => x"a4ec0806",
   578 => x"05795553",
   579 => x"545497d2",
   580 => x"2d029005",
   581 => x"0d04a4f0",
   582 => x"08a0c00c",
   583 => x"0402f405",
   584 => x"0dd45281",
   585 => x"ff720c71",
   586 => x"085381ff",
   587 => x"720c7288",
   588 => x"2b83fe80",
   589 => x"06720870",
   590 => x"81ff0651",
   591 => x"525381ff",
   592 => x"720c7271",
   593 => x"07882b72",
   594 => x"087081ff",
   595 => x"06515253",
   596 => x"81ff720c",
   597 => x"72710788",
   598 => x"2b720870",
   599 => x"81ff0672",
   600 => x"07a0c00c",
   601 => x"5253028c",
   602 => x"050d0402",
   603 => x"f4050d74",
   604 => x"767181ff",
   605 => x"06d40c53",
   606 => x"53a59808",
   607 => x"85387189",
   608 => x"2b527198",
   609 => x"2ad40c71",
   610 => x"902a7081",
   611 => x"ff06d40c",
   612 => x"5171882a",
   613 => x"7081ff06",
   614 => x"d40c5171",
   615 => x"81ff06d4",
   616 => x"0c72902a",
   617 => x"7081ff06",
   618 => x"d40c51d4",
   619 => x"087081ff",
   620 => x"06515182",
   621 => x"b8bf5270",
   622 => x"81ff2e09",
   623 => x"81069438",
   624 => x"81ff0bd4",
   625 => x"0cd40870",
   626 => x"81ff06ff",
   627 => x"14545151",
   628 => x"71e53870",
   629 => x"a0c00c02",
   630 => x"8c050d04",
   631 => x"02fc050d",
   632 => x"81c75181",
   633 => x"ff0bd40c",
   634 => x"ff115170",
   635 => x"8025f438",
   636 => x"0284050d",
   637 => x"0402f005",
   638 => x"0d93dc2d",
   639 => x"8fcf5380",
   640 => x"5287fc80",
   641 => x"f75192eb",
   642 => x"2da0c008",
   643 => x"54a0c008",
   644 => x"812e0981",
   645 => x"06a33881",
   646 => x"ff0bd40c",
   647 => x"820a5284",
   648 => x"9c80e951",
   649 => x"92eb2da0",
   650 => x"c0088b38",
   651 => x"81ff0bd4",
   652 => x"0c735394",
   653 => x"bf0493dc",
   654 => x"2dff1353",
   655 => x"72c13872",
   656 => x"a0c00c02",
   657 => x"90050d04",
   658 => x"02f4050d",
   659 => x"81ff0bd4",
   660 => x"0c935380",
   661 => x"5287fc80",
   662 => x"c15192eb",
   663 => x"2da0c008",
   664 => x"8b3881ff",
   665 => x"0bd40c81",
   666 => x"5394f504",
   667 => x"93dc2dff",
   668 => x"135372df",
   669 => x"3872a0c0",
   670 => x"0c028c05",
   671 => x"0d0402f0",
   672 => x"050d93dc",
   673 => x"2d83aa52",
   674 => x"849c80c8",
   675 => x"5192eb2d",
   676 => x"a0c00881",
   677 => x"2e098106",
   678 => x"9238929d",
   679 => x"2da0c008",
   680 => x"83ffff06",
   681 => x"537283aa",
   682 => x"2e973894",
   683 => x"c82d95bc",
   684 => x"04815496",
   685 => x"a1049fac",
   686 => x"5185f32d",
   687 => x"805496a1",
   688 => x"0481ff0b",
   689 => x"d40cb153",
   690 => x"93f52da0",
   691 => x"c008802e",
   692 => x"80c03880",
   693 => x"5287fc80",
   694 => x"fa5192eb",
   695 => x"2da0c008",
   696 => x"b13881ff",
   697 => x"0bd40cd4",
   698 => x"085381ff",
   699 => x"0bd40c81",
   700 => x"ff0bd40c",
   701 => x"81ff0bd4",
   702 => x"0c81ff0b",
   703 => x"d40c7286",
   704 => x"2a708106",
   705 => x"a0c00856",
   706 => x"51537280",
   707 => x"2e933895",
   708 => x"b1047282",
   709 => x"2eff9f38",
   710 => x"ff135372",
   711 => x"ffaa3872",
   712 => x"5473a0c0",
   713 => x"0c029005",
   714 => x"0d0402f0",
   715 => x"050d810b",
   716 => x"a5980c84",
   717 => x"54d00870",
   718 => x"8f2a7081",
   719 => x"06515153",
   720 => x"72f33872",
   721 => x"d00c93dc",
   722 => x"2d9fbc51",
   723 => x"85f32dd0",
   724 => x"08708f2a",
   725 => x"70810651",
   726 => x"515372f3",
   727 => x"38810bd0",
   728 => x"0cb15380",
   729 => x"5284d480",
   730 => x"c05192eb",
   731 => x"2da0c008",
   732 => x"812ea138",
   733 => x"72822e09",
   734 => x"81068c38",
   735 => x"9fc85185",
   736 => x"f32d8053",
   737 => x"97c904ff",
   738 => x"135372d7",
   739 => x"38ff1454",
   740 => x"73ffa238",
   741 => x"94fe2da0",
   742 => x"c008a598",
   743 => x"0ca0c008",
   744 => x"8b388152",
   745 => x"87fc80d0",
   746 => x"5192eb2d",
   747 => x"81ff0bd4",
   748 => x"0cd00870",
   749 => x"8f2a7081",
   750 => x"06515153",
   751 => x"72f33872",
   752 => x"d00c81ff",
   753 => x"0bd40c81",
   754 => x"5372a0c0",
   755 => x"0c029005",
   756 => x"0d0402e8",
   757 => x"050d7855",
   758 => x"805681ff",
   759 => x"0bd40cd0",
   760 => x"08708f2a",
   761 => x"70810651",
   762 => x"515372f3",
   763 => x"3882810b",
   764 => x"d00c81ff",
   765 => x"0bd40c77",
   766 => x"5287fc80",
   767 => x"d15192eb",
   768 => x"2d80dbc6",
   769 => x"df54a0c0",
   770 => x"08802e8a",
   771 => x"389eac51",
   772 => x"85f32d98",
   773 => x"e40481ff",
   774 => x"0bd40cd4",
   775 => x"087081ff",
   776 => x"06515372",
   777 => x"81fe2e09",
   778 => x"81069d38",
   779 => x"80ff5392",
   780 => x"9d2da0c0",
   781 => x"08757084",
   782 => x"05570cff",
   783 => x"13537280",
   784 => x"25ed3881",
   785 => x"5698ce04",
   786 => x"ff145473",
   787 => x"c93881ff",
   788 => x"0bd40cd0",
   789 => x"08708f2a",
   790 => x"70810651",
   791 => x"515372f3",
   792 => x"3872d00c",
   793 => x"75a0c00c",
   794 => x"0298050d",
   795 => x"04a59808",
   796 => x"a0c00c04",
   797 => x"02f4050d",
   798 => x"7470882a",
   799 => x"83fe8006",
   800 => x"7072982a",
   801 => x"0772882b",
   802 => x"87fc8080",
   803 => x"0673982b",
   804 => x"81f00a06",
   805 => x"71730707",
   806 => x"a0c00c56",
   807 => x"51535102",
   808 => x"8c050d04",
   809 => x"02f8050d",
   810 => x"028e0580",
   811 => x"f52d7488",
   812 => x"2b077083",
   813 => x"ffff06a0",
   814 => x"c00c5102",
   815 => x"88050d04",
   816 => x"02fc050d",
   817 => x"72518071",
   818 => x"0c800b84",
   819 => x"120c0284",
   820 => x"050d0402",
   821 => x"f4050d9d",
   822 => x"a32de008",
   823 => x"e408718b",
   824 => x"2a708106",
   825 => x"51535452",
   826 => x"70802e9d",
   827 => x"38a59c08",
   828 => x"708429a5",
   829 => x"a4057381",
   830 => x"ff06710c",
   831 => x"5151a59c",
   832 => x"08811187",
   833 => x"06a59c0c",
   834 => x"51728b2a",
   835 => x"70810651",
   836 => x"5170802e",
   837 => x"8192389f",
   838 => x"fc088429",
   839 => x"a5d00573",
   840 => x"81ff0671",
   841 => x"0c519ffc",
   842 => x"0881059f",
   843 => x"fc0c850b",
   844 => x"9ff80c9f",
   845 => x"fc089ff4",
   846 => x"082e0981",
   847 => x"0681a638",
   848 => x"800b9ffc",
   849 => x"0ca5e008",
   850 => x"819b38a5",
   851 => x"d0087009",
   852 => x"708306fe",
   853 => x"cc0c5270",
   854 => x"852a7081",
   855 => x"06a5c808",
   856 => x"55515253",
   857 => x"70802e8e",
   858 => x"38a5d808",
   859 => x"fe803212",
   860 => x"a5c80c9a",
   861 => x"fd04a5d8",
   862 => x"0812a5c8",
   863 => x"0c72842a",
   864 => x"708106a5",
   865 => x"c4085451",
   866 => x"5170802e",
   867 => x"9038a5d4",
   868 => x"0881ff32",
   869 => x"128105a5",
   870 => x"c40c9be5",
   871 => x"0471a5d4",
   872 => x"0831a5c4",
   873 => x"0c9be504",
   874 => x"9ff808ff",
   875 => x"059ff80c",
   876 => x"9ff808ff",
   877 => x"2e098106",
   878 => x"ac389ffc",
   879 => x"08802e92",
   880 => x"38810ba5",
   881 => x"e00c870b",
   882 => x"9ff40831",
   883 => x"9ff40c9b",
   884 => x"e004a5e0",
   885 => x"08517080",
   886 => x"2e8638ff",
   887 => x"11a5e00c",
   888 => x"800b9ffc",
   889 => x"0c800ba5",
   890 => x"cc0c9d96",
   891 => x"2d9d9d2d",
   892 => x"028c050d",
   893 => x"0402fc05",
   894 => x"0d9da32d",
   895 => x"810ba5cc",
   896 => x"0c9d9d2d",
   897 => x"a5cc0851",
   898 => x"70fa3802",
   899 => x"84050d04",
   900 => x"02f8050d",
   901 => x"a59c5199",
   902 => x"c02d800b",
   903 => x"a5e00c83",
   904 => x"0b9ff40c",
   905 => x"e408708c",
   906 => x"2a708106",
   907 => x"51515271",
   908 => x"802e8638",
   909 => x"840b9ff4",
   910 => x"0ce40870",
   911 => x"8d2a7081",
   912 => x"06515152",
   913 => x"71802e9f",
   914 => x"38870b9f",
   915 => x"f408319f",
   916 => x"f40ce408",
   917 => x"708a2a70",
   918 => x"81065151",
   919 => x"5271802e",
   920 => x"f13881f4",
   921 => x"0be40c99",
   922 => x"d3519d92",
   923 => x"2d9cf52d",
   924 => x"0288050d",
   925 => x"0402f805",
   926 => x"0da08052",
   927 => x"8f518072",
   928 => x"70840554",
   929 => x"0cff1151",
   930 => x"708025f2",
   931 => x"38028805",
   932 => x"0d047198",
   933 => x"0c04ffb0",
   934 => x"08a0c00c",
   935 => x"04810bff",
   936 => x"b00c0480",
   937 => x"0bffb00c",
   938 => x"04000000",
   939 => x"00ffffff",
   940 => x"ff00ffff",
   941 => x"ffff00ff",
   942 => x"ffffff00",
   943 => x"496e6974",
   944 => x"69616c69",
   945 => x"7a696e67",
   946 => x"20534420",
   947 => x"63617264",
   948 => x"0a000000",
   949 => x"53444843",
   950 => x"20636172",
   951 => x"64206465",
   952 => x"74656374",
   953 => x"65640a00",
   954 => x"46617433",
   955 => x"32206465",
   956 => x"74656374",
   957 => x"65640a00",
   958 => x"54727969",
   959 => x"6e672053",
   960 => x"50454343",
   961 => x"592e524f",
   962 => x"4d0a0000",
   963 => x"53504543",
   964 => x"43592020",
   965 => x"524f4d00",
   966 => x"4c6f6164",
   967 => x"696e6720",
   968 => x"53504543",
   969 => x"43592e52",
   970 => x"4f4d0a00",
   971 => x"52656164",
   972 => x"20666169",
   973 => x"6c65640a",
   974 => x"00000000",
   975 => x"4c6f6164",
   976 => x"696e6720",
   977 => x"42494f53",
   978 => x"20646f6e",
   979 => x"650a0000",
   980 => x"4c6f6164",
   981 => x"696e6720",
   982 => x"42494f53",
   983 => x"20666169",
   984 => x"6c65640a",
   985 => x"00000000",
   986 => x"4d425220",
   987 => x"6661696c",
   988 => x"0a000000",
   989 => x"46415431",
   990 => x"36202020",
   991 => x"00000000",
   992 => x"46415433",
   993 => x"32202020",
   994 => x"00000000",
   995 => x"4e6f2070",
   996 => x"61727469",
   997 => x"74696f6e",
   998 => x"20736967",
   999 => x"0a000000",
  1000 => x"42616420",
  1001 => x"70617274",
  1002 => x"0a000000",
  1003 => x"53444843",
  1004 => x"20657272",
  1005 => x"6f72210a",
  1006 => x"00000000",
  1007 => x"53442069",
  1008 => x"6e69742e",
  1009 => x"2e2e0a00",
  1010 => x"53442063",
  1011 => x"61726420",
  1012 => x"72657365",
  1013 => x"74206661",
  1014 => x"696c6564",
  1015 => x"210a0000",
  1016 => x"57726974",
  1017 => x"65206661",
  1018 => x"696c6564",
  1019 => x"0a000000",
  1020 => x"00000002",
  1021 => x"00000003",
  1022 => x"00000000",
  1023 => x"00000000",
  1024 => x"00000000",
  1025 => x"00000000",
  1026 => x"00000000",
  1027 => x"00000000",
  1028 => x"00000000",
  1029 => x"00000000",
  1030 => x"00000000",
  1031 => x"00000000",
  1032 => x"00000000",
  1033 => x"00000000",
  1034 => x"00000000",
  1035 => x"00000000",
  1036 => x"00000000",
  1037 => x"00000000",
  1038 => x"00000000",
  1039 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

