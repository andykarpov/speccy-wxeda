-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity loader_firmware_rom is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end loader_firmware_rom;

architecture arch of loader_firmware_rom is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0ba9",
     9 => x"d8080b0b",
    10 => x"0ba9dc08",
    11 => x"0b0b0ba9",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"a9e00c0b",
    16 => x"0b0ba9dc",
    17 => x"0c0b0b0b",
    18 => x"a9d80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba0fc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"a9d870af",
    57 => x"8c278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"89d00402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"a9e80c9f",
    65 => x"0ba9ec0c",
    66 => x"a0717081",
    67 => x"055334a9",
    68 => x"ec08ff05",
    69 => x"a9ec0ca9",
    70 => x"ec088025",
    71 => x"eb38a9e8",
    72 => x"08ff05a9",
    73 => x"e80ca9e8",
    74 => x"088025d7",
    75 => x"38028405",
    76 => x"0d0402f0",
    77 => x"050df880",
    78 => x"53f8a054",
    79 => x"83bf5273",
    80 => x"70810555",
    81 => x"33517073",
    82 => x"70810555",
    83 => x"34ff1252",
    84 => x"718025eb",
    85 => x"38fbc053",
    86 => x"9f52a073",
    87 => x"70810555",
    88 => x"34ff1252",
    89 => x"718025f2",
    90 => x"38029005",
    91 => x"0d0402f4",
    92 => x"050d7453",
    93 => x"8e0ba9e8",
    94 => x"08258f38",
    95 => x"82b22da9",
    96 => x"e808ff05",
    97 => x"a9e80c82",
    98 => x"f404a9e8",
    99 => x"08a9ec08",
   100 => x"5351728a",
   101 => x"2e098106",
   102 => x"b7387151",
   103 => x"719f24a0",
   104 => x"38a9e808",
   105 => x"a02911f8",
   106 => x"80115151",
   107 => x"a07134a9",
   108 => x"ec088105",
   109 => x"a9ec0ca9",
   110 => x"ec08519f",
   111 => x"7125e238",
   112 => x"800ba9ec",
   113 => x"0ca9e808",
   114 => x"8105a9e8",
   115 => x"0c83e404",
   116 => x"70a02912",
   117 => x"f8801151",
   118 => x"51727134",
   119 => x"a9ec0881",
   120 => x"05a9ec0c",
   121 => x"a9ec08a0",
   122 => x"2e098106",
   123 => x"8e38800b",
   124 => x"a9ec0ca9",
   125 => x"e8088105",
   126 => x"a9e80c02",
   127 => x"8c050d04",
   128 => x"02e8050d",
   129 => x"77795656",
   130 => x"880bfc16",
   131 => x"77712c8f",
   132 => x"06545254",
   133 => x"80537272",
   134 => x"25953871",
   135 => x"53fbe014",
   136 => x"51877134",
   137 => x"8114ff14",
   138 => x"545472f1",
   139 => x"387153f9",
   140 => x"1576712c",
   141 => x"87065351",
   142 => x"71802e8b",
   143 => x"38fbe014",
   144 => x"51717134",
   145 => x"81145472",
   146 => x"8e249538",
   147 => x"8f733153",
   148 => x"fbe01451",
   149 => x"a0713481",
   150 => x"14ff1454",
   151 => x"5472f138",
   152 => x"0298050d",
   153 => x"0402ec05",
   154 => x"0d800ba9",
   155 => x"f00cf68c",
   156 => x"08f69008",
   157 => x"71882c56",
   158 => x"5481ff06",
   159 => x"52737225",
   160 => x"88387154",
   161 => x"820ba9f0",
   162 => x"0c72882c",
   163 => x"7381ff06",
   164 => x"54557473",
   165 => x"258b3872",
   166 => x"a9f00884",
   167 => x"07a9f00c",
   168 => x"5573842b",
   169 => x"86a07125",
   170 => x"83713170",
   171 => x"0b0b0ba6",
   172 => x"c00c8171",
   173 => x"2bff05f6",
   174 => x"880cfecc",
   175 => x"13ff122c",
   176 => x"788829ff",
   177 => x"94057081",
   178 => x"2ca9f008",
   179 => x"52585255",
   180 => x"51525476",
   181 => x"802e8538",
   182 => x"70810751",
   183 => x"70f6940c",
   184 => x"71098105",
   185 => x"f6800c72",
   186 => x"098105f6",
   187 => x"840c0294",
   188 => x"050d0402",
   189 => x"f4050d74",
   190 => x"53727081",
   191 => x"055480f5",
   192 => x"2d527180",
   193 => x"2e893871",
   194 => x"5182ee2d",
   195 => x"85f90402",
   196 => x"8c050d04",
   197 => x"02d4050d",
   198 => x"a3fc5185",
   199 => x"f32d988c",
   200 => x"2da9d808",
   201 => x"802e81ef",
   202 => x"388afb2d",
   203 => x"a9d80853",
   204 => x"a9d80880",
   205 => x"2e81e238",
   206 => x"9acf2da9",
   207 => x"d808802e",
   208 => x"8738a494",
   209 => x"5186d504",
   210 => x"93f82da9",
   211 => x"d808802e",
   212 => x"8738a4a8",
   213 => x"5185f32d",
   214 => x"a4c05185",
   215 => x"f32da4d4",
   216 => x"52a9f451",
   217 => x"918d2da9",
   218 => x"d808802e",
   219 => x"81a938a4",
   220 => x"e05185f3",
   221 => x"2da9f808",
   222 => x"57807759",
   223 => x"5a767a2e",
   224 => x"8b38811a",
   225 => x"78812a59",
   226 => x"5a77f738",
   227 => x"f71a5a80",
   228 => x"772580fe",
   229 => x"38795277",
   230 => x"5184802d",
   231 => x"aa8052a9",
   232 => x"f45193d2",
   233 => x"2da9d808",
   234 => x"53a9d808",
   235 => x"802e80c9",
   236 => x"38aa805b",
   237 => x"805987e6",
   238 => x"047a7084",
   239 => x"055c0870",
   240 => x"81ff0671",
   241 => x"882c7081",
   242 => x"ff067390",
   243 => x"2c7081ff",
   244 => x"0675982a",
   245 => x"fec80cfe",
   246 => x"c80c58fe",
   247 => x"c80c57fe",
   248 => x"c80c841a",
   249 => x"5a537653",
   250 => x"84807725",
   251 => x"84388480",
   252 => x"53727924",
   253 => x"c4388882",
   254 => x"04a4f051",
   255 => x"85f32d88",
   256 => x"9904a9f4",
   257 => x"5193a52d",
   258 => x"fc801781",
   259 => x"19595787",
   260 => x"8f048153",
   261 => x"88990480",
   262 => x"5372a9d8",
   263 => x"0c02ac05",
   264 => x"0d0402f8",
   265 => x"050d9f8b",
   266 => x"2d81f72d",
   267 => x"815184e5",
   268 => x"2dfec452",
   269 => x"81720c9d",
   270 => x"d72d9dd7",
   271 => x"2d84720c",
   272 => x"73518694",
   273 => x"2da78c51",
   274 => x"a0e92d80",
   275 => x"5184e52d",
   276 => x"0288050d",
   277 => x"0402fc05",
   278 => x"0d825188",
   279 => x"a22d0284",
   280 => x"050d0402",
   281 => x"fc050d80",
   282 => x"5188a22d",
   283 => x"0284050d",
   284 => x"0402f405",
   285 => x"0d747081",
   286 => x"8432aefc",
   287 => x"0c708306",
   288 => x"525370a7",
   289 => x"ec0b8805",
   290 => x"81b72d72",
   291 => x"892a7081",
   292 => x"06515170",
   293 => x"a8bc0b81",
   294 => x"b72d7283",
   295 => x"2a810673",
   296 => x"882a7081",
   297 => x"06515252",
   298 => x"70802e85",
   299 => x"38718207",
   300 => x"5271a898",
   301 => x"0b81b72d",
   302 => x"72842c70",
   303 => x"83065151",
   304 => x"70a8a40b",
   305 => x"81b72d70",
   306 => x"a9d80c02",
   307 => x"8c050d04",
   308 => x"02f8050d",
   309 => x"84b85188",
   310 => x"f12d810b",
   311 => x"fec40c84",
   312 => x"b80bfec0",
   313 => x"0c840bfe",
   314 => x"c40c830b",
   315 => x"fecc0c9d",
   316 => x"f22d9eff",
   317 => x"2d9dd72d",
   318 => x"9dd72d81",
   319 => x"f72d8151",
   320 => x"84e52d9d",
   321 => x"d72d9dd7",
   322 => x"2d80ff52",
   323 => x"9dd72d81",
   324 => x"5184e52d",
   325 => x"ff125271",
   326 => x"8025f138",
   327 => x"9dd72d9d",
   328 => x"d72d8151",
   329 => x"86942da9",
   330 => x"d808802e",
   331 => x"8738a580",
   332 => x"518ab704",
   333 => x"a5945185",
   334 => x"f32d8aa2",
   335 => x"0402e805",
   336 => x"0d77797b",
   337 => x"58555580",
   338 => x"53727625",
   339 => x"a3387470",
   340 => x"81055680",
   341 => x"f52d7470",
   342 => x"81055680",
   343 => x"f52d5252",
   344 => x"71712e86",
   345 => x"3881518a",
   346 => x"f2048113",
   347 => x"538ac904",
   348 => x"805170a9",
   349 => x"d80c0298",
   350 => x"050d0402",
   351 => x"d8050d80",
   352 => x"0bae880c",
   353 => x"aa805280",
   354 => x"5199b42d",
   355 => x"a9d80854",
   356 => x"a9d8088c",
   357 => x"38a5ac51",
   358 => x"85f32d73",
   359 => x"55909604",
   360 => x"8056810b",
   361 => x"aeac0c88",
   362 => x"53a5b852",
   363 => x"aab6518a",
   364 => x"bd2da9d8",
   365 => x"08762e09",
   366 => x"81068738",
   367 => x"a9d808ae",
   368 => x"ac0c8853",
   369 => x"a5c452aa",
   370 => x"d2518abd",
   371 => x"2da9d808",
   372 => x"8738a9d8",
   373 => x"08aeac0c",
   374 => x"aeac0880",
   375 => x"2e80f638",
   376 => x"adc60b80",
   377 => x"f52dadc7",
   378 => x"0b80f52d",
   379 => x"71982b71",
   380 => x"902b07ad",
   381 => x"c80b80f5",
   382 => x"2d70882b",
   383 => x"7207adc9",
   384 => x"0b80f52d",
   385 => x"7107adfe",
   386 => x"0b80f52d",
   387 => x"adff0b80",
   388 => x"f52d7188",
   389 => x"2b07535f",
   390 => x"54525a56",
   391 => x"57557381",
   392 => x"abaa2e09",
   393 => x"81068d38",
   394 => x"75519ad6",
   395 => x"2da9d808",
   396 => x"568cc104",
   397 => x"7382d4d5",
   398 => x"2e8738a5",
   399 => x"d0518d82",
   400 => x"04aa8052",
   401 => x"755199b4",
   402 => x"2da9d808",
   403 => x"55a9d808",
   404 => x"802e83c2",
   405 => x"388853a5",
   406 => x"c452aad2",
   407 => x"518abd2d",
   408 => x"a9d80889",
   409 => x"38810bae",
   410 => x"880c8d88",
   411 => x"048853a5",
   412 => x"b852aab6",
   413 => x"518abd2d",
   414 => x"a9d80880",
   415 => x"2e8a38a5",
   416 => x"e45185f3",
   417 => x"2d8de204",
   418 => x"adfe0b80",
   419 => x"f52d5473",
   420 => x"80d52e09",
   421 => x"810680ca",
   422 => x"38adff0b",
   423 => x"80f52d54",
   424 => x"7381aa2e",
   425 => x"098106ba",
   426 => x"38800baa",
   427 => x"800b80f5",
   428 => x"2d565474",
   429 => x"81e92e83",
   430 => x"38815474",
   431 => x"81eb2e8c",
   432 => x"38805573",
   433 => x"752e0981",
   434 => x"0682cb38",
   435 => x"aa8b0b80",
   436 => x"f52d5574",
   437 => x"8d38aa8c",
   438 => x"0b80f52d",
   439 => x"5473822e",
   440 => x"86388055",
   441 => x"909604aa",
   442 => x"8d0b80f5",
   443 => x"2d70ae80",
   444 => x"0cff05ae",
   445 => x"840caa8e",
   446 => x"0b80f52d",
   447 => x"aa8f0b80",
   448 => x"f52d5876",
   449 => x"05778280",
   450 => x"290570ae",
   451 => x"8c0caa90",
   452 => x"0b80f52d",
   453 => x"70aea00c",
   454 => x"ae880859",
   455 => x"57587680",
   456 => x"2e81a338",
   457 => x"8853a5c4",
   458 => x"52aad251",
   459 => x"8abd2da9",
   460 => x"d80881e2",
   461 => x"38ae8008",
   462 => x"70842bae",
   463 => x"a40c70ae",
   464 => x"9c0caaa5",
   465 => x"0b80f52d",
   466 => x"aaa40b80",
   467 => x"f52d7182",
   468 => x"802905aa",
   469 => x"a60b80f5",
   470 => x"2d708480",
   471 => x"802912aa",
   472 => x"a70b80f5",
   473 => x"2d708180",
   474 => x"0a291270",
   475 => x"aea80cae",
   476 => x"a0087129",
   477 => x"ae8c0805",
   478 => x"70ae900c",
   479 => x"aaad0b80",
   480 => x"f52daaac",
   481 => x"0b80f52d",
   482 => x"71828029",
   483 => x"05aaae0b",
   484 => x"80f52d70",
   485 => x"84808029",
   486 => x"12aaaf0b",
   487 => x"80f52d70",
   488 => x"982b81f0",
   489 => x"0a067205",
   490 => x"70ae940c",
   491 => x"fe117e29",
   492 => x"7705ae98",
   493 => x"0c525952",
   494 => x"43545e51",
   495 => x"5259525d",
   496 => x"57595790",
   497 => x"9404aa92",
   498 => x"0b80f52d",
   499 => x"aa910b80",
   500 => x"f52d7182",
   501 => x"80290570",
   502 => x"aea40c70",
   503 => x"a02983ff",
   504 => x"0570892a",
   505 => x"70ae9c0c",
   506 => x"aa970b80",
   507 => x"f52daa96",
   508 => x"0b80f52d",
   509 => x"71828029",
   510 => x"0570aea8",
   511 => x"0c7b7129",
   512 => x"1e70ae98",
   513 => x"0c7dae94",
   514 => x"0c7305ae",
   515 => x"900c555e",
   516 => x"51515555",
   517 => x"815574a9",
   518 => x"d80c02a8",
   519 => x"050d0402",
   520 => x"ec050d76",
   521 => x"70872c71",
   522 => x"80ff0655",
   523 => x"5654ae88",
   524 => x"088a3873",
   525 => x"882c7481",
   526 => x"ff065455",
   527 => x"aa8052ae",
   528 => x"8c081551",
   529 => x"99b42da9",
   530 => x"d80854a9",
   531 => x"d808802e",
   532 => x"b338ae88",
   533 => x"08802e98",
   534 => x"38728429",
   535 => x"aa800570",
   536 => x"0852539a",
   537 => x"d62da9d8",
   538 => x"08f00a06",
   539 => x"53918204",
   540 => x"7210aa80",
   541 => x"057080e0",
   542 => x"2d52539b",
   543 => x"862da9d8",
   544 => x"08537254",
   545 => x"73a9d80c",
   546 => x"0294050d",
   547 => x"0402c805",
   548 => x"0d7f615f",
   549 => x"5b800bae",
   550 => x"9408ae98",
   551 => x"08595d56",
   552 => x"ae880876",
   553 => x"2e8a38ae",
   554 => x"8008842b",
   555 => x"5891b604",
   556 => x"ae9c0884",
   557 => x"2b588059",
   558 => x"78782781",
   559 => x"a938788f",
   560 => x"06a01757",
   561 => x"54738f38",
   562 => x"aa805276",
   563 => x"51811757",
   564 => x"99b42daa",
   565 => x"80568076",
   566 => x"80f52d56",
   567 => x"5474742e",
   568 => x"83388154",
   569 => x"7481e52e",
   570 => x"80f63881",
   571 => x"70750655",
   572 => x"5d73802e",
   573 => x"80ea388b",
   574 => x"1680f52d",
   575 => x"98065a79",
   576 => x"80de388b",
   577 => x"537d5275",
   578 => x"518abd2d",
   579 => x"a9d80880",
   580 => x"cf389c16",
   581 => x"08519ad6",
   582 => x"2da9d808",
   583 => x"841c0c9a",
   584 => x"1680e02d",
   585 => x"519b862d",
   586 => x"a9d808a9",
   587 => x"d808881d",
   588 => x"0ca9d808",
   589 => x"5555ae88",
   590 => x"08802e98",
   591 => x"38941680",
   592 => x"e02d519b",
   593 => x"862da9d8",
   594 => x"08902b83",
   595 => x"fff00a06",
   596 => x"70165154",
   597 => x"73881c0c",
   598 => x"797b0c7c",
   599 => x"54939c04",
   600 => x"81195991",
   601 => x"b804ae88",
   602 => x"08802eae",
   603 => x"387b5190",
   604 => x"9f2da9d8",
   605 => x"08a9d808",
   606 => x"80ffffff",
   607 => x"f806555c",
   608 => x"7380ffff",
   609 => x"fff82e92",
   610 => x"38a9d808",
   611 => x"fe05ae80",
   612 => x"0829ae90",
   613 => x"08055791",
   614 => x"b6048054",
   615 => x"73a9d80c",
   616 => x"02b8050d",
   617 => x"0402f405",
   618 => x"0d747008",
   619 => x"8105710c",
   620 => x"7008ae84",
   621 => x"08065353",
   622 => x"718e3888",
   623 => x"13085190",
   624 => x"9f2da9d8",
   625 => x"0888140c",
   626 => x"810ba9d8",
   627 => x"0c028c05",
   628 => x"0d0402f0",
   629 => x"050d7588",
   630 => x"1108fe05",
   631 => x"ae800829",
   632 => x"ae900811",
   633 => x"7208ae84",
   634 => x"08060579",
   635 => x"55535454",
   636 => x"99b42d02",
   637 => x"90050d04",
   638 => x"ae8808a9",
   639 => x"d80c0402",
   640 => x"f4050dd4",
   641 => x"5281ff72",
   642 => x"0c710853",
   643 => x"81ff720c",
   644 => x"72882b83",
   645 => x"fe800672",
   646 => x"087081ff",
   647 => x"06515253",
   648 => x"81ff720c",
   649 => x"72710788",
   650 => x"2b720870",
   651 => x"81ff0651",
   652 => x"525381ff",
   653 => x"720c7271",
   654 => x"07882b72",
   655 => x"087081ff",
   656 => x"067207a9",
   657 => x"d80c5253",
   658 => x"028c050d",
   659 => x"0402f405",
   660 => x"0d747671",
   661 => x"81ff06d4",
   662 => x"0c5353ae",
   663 => x"b0088538",
   664 => x"71892b52",
   665 => x"71982ad4",
   666 => x"0c71902a",
   667 => x"7081ff06",
   668 => x"d40c5171",
   669 => x"882a7081",
   670 => x"ff06d40c",
   671 => x"517181ff",
   672 => x"06d40c72",
   673 => x"902a7081",
   674 => x"ff06d40c",
   675 => x"51d40870",
   676 => x"81ff0651",
   677 => x"5182b8bf",
   678 => x"527081ff",
   679 => x"2e098106",
   680 => x"943881ff",
   681 => x"0bd40cd4",
   682 => x"087081ff",
   683 => x"06ff1454",
   684 => x"515171e5",
   685 => x"3870a9d8",
   686 => x"0c028c05",
   687 => x"0d0402fc",
   688 => x"050d81c7",
   689 => x"5181ff0b",
   690 => x"d40cff11",
   691 => x"51708025",
   692 => x"f4380284",
   693 => x"050d0402",
   694 => x"f0050d95",
   695 => x"be2d8fcf",
   696 => x"53805287",
   697 => x"fc80f751",
   698 => x"94cd2da9",
   699 => x"d80854a9",
   700 => x"d808812e",
   701 => x"098106a3",
   702 => x"3881ff0b",
   703 => x"d40c820a",
   704 => x"52849c80",
   705 => x"e95194cd",
   706 => x"2da9d808",
   707 => x"8b3881ff",
   708 => x"0bd40c73",
   709 => x"5396a104",
   710 => x"95be2dff",
   711 => x"135372c1",
   712 => x"3872a9d8",
   713 => x"0c029005",
   714 => x"0d0402f4",
   715 => x"050d81ff",
   716 => x"0bd40c93",
   717 => x"53805287",
   718 => x"fc80c151",
   719 => x"94cd2da9",
   720 => x"d8088b38",
   721 => x"81ff0bd4",
   722 => x"0c815396",
   723 => x"d70495be",
   724 => x"2dff1353",
   725 => x"72df3872",
   726 => x"a9d80c02",
   727 => x"8c050d04",
   728 => x"02f0050d",
   729 => x"95be2d83",
   730 => x"aa52849c",
   731 => x"80c85194",
   732 => x"cd2da9d8",
   733 => x"08812e09",
   734 => x"81069238",
   735 => x"93ff2da9",
   736 => x"d80883ff",
   737 => x"ff065372",
   738 => x"83aa2e97",
   739 => x"3896aa2d",
   740 => x"979e0481",
   741 => x"54988304",
   742 => x"a5f05185",
   743 => x"f32d8054",
   744 => x"98830481",
   745 => x"ff0bd40c",
   746 => x"b15395d7",
   747 => x"2da9d808",
   748 => x"802e80c0",
   749 => x"38805287",
   750 => x"fc80fa51",
   751 => x"94cd2da9",
   752 => x"d808b138",
   753 => x"81ff0bd4",
   754 => x"0cd40853",
   755 => x"81ff0bd4",
   756 => x"0c81ff0b",
   757 => x"d40c81ff",
   758 => x"0bd40c81",
   759 => x"ff0bd40c",
   760 => x"72862a70",
   761 => x"8106a9d8",
   762 => x"08565153",
   763 => x"72802e93",
   764 => x"38979304",
   765 => x"72822eff",
   766 => x"9f38ff13",
   767 => x"5372ffaa",
   768 => x"38725473",
   769 => x"a9d80c02",
   770 => x"90050d04",
   771 => x"02f0050d",
   772 => x"810baeb0",
   773 => x"0c8454d0",
   774 => x"08708f2a",
   775 => x"70810651",
   776 => x"515372f3",
   777 => x"3872d00c",
   778 => x"95be2da6",
   779 => x"805185f3",
   780 => x"2dd00870",
   781 => x"8f2a7081",
   782 => x"06515153",
   783 => x"72f33881",
   784 => x"0bd00cb1",
   785 => x"53805284",
   786 => x"d480c051",
   787 => x"94cd2da9",
   788 => x"d808812e",
   789 => x"a1387282",
   790 => x"2e098106",
   791 => x"8c38a68c",
   792 => x"5185f32d",
   793 => x"805399ab",
   794 => x"04ff1353",
   795 => x"72d738ff",
   796 => x"145473ff",
   797 => x"a23896e0",
   798 => x"2da9d808",
   799 => x"aeb00ca9",
   800 => x"d8088b38",
   801 => x"815287fc",
   802 => x"80d05194",
   803 => x"cd2d81ff",
   804 => x"0bd40cd0",
   805 => x"08708f2a",
   806 => x"70810651",
   807 => x"515372f3",
   808 => x"3872d00c",
   809 => x"81ff0bd4",
   810 => x"0c815372",
   811 => x"a9d80c02",
   812 => x"90050d04",
   813 => x"02e8050d",
   814 => x"78558056",
   815 => x"81ff0bd4",
   816 => x"0cd00870",
   817 => x"8f2a7081",
   818 => x"06515153",
   819 => x"72f33882",
   820 => x"810bd00c",
   821 => x"81ff0bd4",
   822 => x"0c775287",
   823 => x"fc80d151",
   824 => x"94cd2d80",
   825 => x"dbc6df54",
   826 => x"a9d80880",
   827 => x"2e8a38a4",
   828 => x"f05185f3",
   829 => x"2d9ac604",
   830 => x"81ff0bd4",
   831 => x"0cd40870",
   832 => x"81ff0651",
   833 => x"537281fe",
   834 => x"2e098106",
   835 => x"9d3880ff",
   836 => x"5393ff2d",
   837 => x"a9d80875",
   838 => x"70840557",
   839 => x"0cff1353",
   840 => x"728025ed",
   841 => x"3881569a",
   842 => x"b004ff14",
   843 => x"5473c938",
   844 => x"81ff0bd4",
   845 => x"0cd00870",
   846 => x"8f2a7081",
   847 => x"06515153",
   848 => x"72f33872",
   849 => x"d00c75a9",
   850 => x"d80c0298",
   851 => x"050d04ae",
   852 => x"b008a9d8",
   853 => x"0c0402f4",
   854 => x"050d7470",
   855 => x"882a83fe",
   856 => x"80067072",
   857 => x"982a0772",
   858 => x"882b87fc",
   859 => x"80800673",
   860 => x"982b81f0",
   861 => x"0a067173",
   862 => x"0707a9d8",
   863 => x"0c565153",
   864 => x"51028c05",
   865 => x"0d0402f8",
   866 => x"050d028e",
   867 => x"0580f52d",
   868 => x"74882b07",
   869 => x"7083ffff",
   870 => x"06a9d80c",
   871 => x"51028805",
   872 => x"0d0402fc",
   873 => x"050d7251",
   874 => x"80710c80",
   875 => x"0b84120c",
   876 => x"0284050d",
   877 => x"0402f405",
   878 => x"0d9f852d",
   879 => x"e008e408",
   880 => x"718b2a70",
   881 => x"81065153",
   882 => x"54527080",
   883 => x"2e9d38ae",
   884 => x"b4087084",
   885 => x"29aebc05",
   886 => x"7381ff06",
   887 => x"710c5151",
   888 => x"aeb40881",
   889 => x"118706ae",
   890 => x"b40c5172",
   891 => x"8b2a7081",
   892 => x"06515170",
   893 => x"802e8192",
   894 => x"38a99008",
   895 => x"8429aee8",
   896 => x"057381ff",
   897 => x"06710c51",
   898 => x"a9900881",
   899 => x"05a9900c",
   900 => x"850ba98c",
   901 => x"0ca99008",
   902 => x"a988082e",
   903 => x"09810681",
   904 => x"a638800b",
   905 => x"a9900cae",
   906 => x"f808819b",
   907 => x"38aee808",
   908 => x"70097083",
   909 => x"06fecc0c",
   910 => x"5270852a",
   911 => x"708106ae",
   912 => x"e0085551",
   913 => x"52537080",
   914 => x"2e8e38ae",
   915 => x"f008fe80",
   916 => x"3212aee0",
   917 => x"0c9cdf04",
   918 => x"aef00812",
   919 => x"aee00c72",
   920 => x"842a7081",
   921 => x"06aedc08",
   922 => x"54515170",
   923 => x"802e9038",
   924 => x"aeec0881",
   925 => x"ff321281",
   926 => x"05aedc0c",
   927 => x"9dc70471",
   928 => x"aeec0831",
   929 => x"aedc0c9d",
   930 => x"c704a98c",
   931 => x"08ff05a9",
   932 => x"8c0ca98c",
   933 => x"08ff2e09",
   934 => x"8106ac38",
   935 => x"a9900880",
   936 => x"2e923881",
   937 => x"0baef80c",
   938 => x"870ba988",
   939 => x"0831a988",
   940 => x"0c9dc204",
   941 => x"aef80851",
   942 => x"70802e86",
   943 => x"38ff11ae",
   944 => x"f80c800b",
   945 => x"a9900c80",
   946 => x"0baee40c",
   947 => x"9ef82d9e",
   948 => x"ff2d028c",
   949 => x"050d0402",
   950 => x"fc050d9f",
   951 => x"852d810b",
   952 => x"aee40c9e",
   953 => x"ff2daee4",
   954 => x"085170fa",
   955 => x"38028405",
   956 => x"0d0402f8",
   957 => x"050daeb4",
   958 => x"519ba22d",
   959 => x"800baef8",
   960 => x"0c830ba9",
   961 => x"880ce408",
   962 => x"708c2a70",
   963 => x"81065151",
   964 => x"5271802e",
   965 => x"8638840b",
   966 => x"a9880ce4",
   967 => x"08708d2a",
   968 => x"70810651",
   969 => x"51527180",
   970 => x"2e9f3887",
   971 => x"0ba98808",
   972 => x"31a9880c",
   973 => x"e408708a",
   974 => x"2a708106",
   975 => x"51515271",
   976 => x"802ef138",
   977 => x"81f40be4",
   978 => x"0c9bb551",
   979 => x"9ef42d9e",
   980 => x"d72d0288",
   981 => x"050d0402",
   982 => x"f8050da9",
   983 => x"94528f51",
   984 => x"80727084",
   985 => x"05540cff",
   986 => x"11517080",
   987 => x"25f23802",
   988 => x"88050d04",
   989 => x"71980c04",
   990 => x"ffb008a9",
   991 => x"d80c0481",
   992 => x"0bffb00c",
   993 => x"04800bff",
   994 => x"b00c0402",
   995 => x"fc050d80",
   996 => x"0ba9d40c",
   997 => x"805184e5",
   998 => x"2d028405",
   999 => x"0d0402ec",
  1000 => x"050d7654",
  1001 => x"8052870b",
  1002 => x"881580f5",
  1003 => x"2d565374",
  1004 => x"72248338",
  1005 => x"a0537251",
  1006 => x"82ee2d81",
  1007 => x"128b1580",
  1008 => x"f52d5452",
  1009 => x"727225de",
  1010 => x"38029405",
  1011 => x"0d0402f0",
  1012 => x"050daf80",
  1013 => x"085481f7",
  1014 => x"2d800baf",
  1015 => x"840c7308",
  1016 => x"802e8180",
  1017 => x"38820ba9",
  1018 => x"ec0caf84",
  1019 => x"088f06a9",
  1020 => x"e80c7308",
  1021 => x"5271832e",
  1022 => x"96387183",
  1023 => x"26893871",
  1024 => x"812eaf38",
  1025 => x"a0cf0471",
  1026 => x"852e9f38",
  1027 => x"a0cf0488",
  1028 => x"1480f52d",
  1029 => x"841508a6",
  1030 => x"b4535452",
  1031 => x"85f32d71",
  1032 => x"84291370",
  1033 => x"085252a0",
  1034 => x"d3047351",
  1035 => x"9f9e2da0",
  1036 => x"cf04aefc",
  1037 => x"08881508",
  1038 => x"2c708106",
  1039 => x"51527180",
  1040 => x"2e8738a6",
  1041 => x"b851a0cc",
  1042 => x"04a6bc51",
  1043 => x"85f32d84",
  1044 => x"14085185",
  1045 => x"f32daf84",
  1046 => x"088105af",
  1047 => x"840c8c14",
  1048 => x"549fde04",
  1049 => x"0290050d",
  1050 => x"0471af80",
  1051 => x"0c9fce2d",
  1052 => x"af8408ff",
  1053 => x"05af880c",
  1054 => x"04000000",
  1055 => x"00ffffff",
  1056 => x"ff00ffff",
  1057 => x"ffff00ff",
  1058 => x"ffffff00",
  1059 => x"4d617374",
  1060 => x"65720000",
  1061 => x"4f504c4c",
  1062 => x"00000000",
  1063 => x"53434300",
  1064 => x"50534700",
  1065 => x"4261636b",
  1066 => x"00000000",
  1067 => x"52657365",
  1068 => x"74000000",
  1069 => x"53617665",
  1070 => x"20616e64",
  1071 => x"20526573",
  1072 => x"65740000",
  1073 => x"4f707469",
  1074 => x"6f6e7320",
  1075 => x"10000000",
  1076 => x"536f756e",
  1077 => x"64201000",
  1078 => x"54757262",
  1079 => x"6f000000",
  1080 => x"4d6f7573",
  1081 => x"6520656d",
  1082 => x"756c6174",
  1083 => x"696f6e00",
  1084 => x"45786974",
  1085 => x"00000000",
  1086 => x"5363616e",
  1087 => x"6c696e65",
  1088 => x"73000000",
  1089 => x"53442043",
  1090 => x"61726400",
  1091 => x"4a617061",
  1092 => x"6e657365",
  1093 => x"206b6579",
  1094 => x"206c6179",
  1095 => x"6f757400",
  1096 => x"32303438",
  1097 => x"4b422052",
  1098 => x"414d0000",
  1099 => x"34303936",
  1100 => x"4b422052",
  1101 => x"414d0000",
  1102 => x"536c323a",
  1103 => x"204e6f6e",
  1104 => x"65000000",
  1105 => x"536c323a",
  1106 => x"20455345",
  1107 => x"2d534343",
  1108 => x"20314d42",
  1109 => x"2f534343",
  1110 => x"2d490000",
  1111 => x"536c323a",
  1112 => x"20455345",
  1113 => x"2d52414d",
  1114 => x"20314d42",
  1115 => x"2f415343",
  1116 => x"49493800",
  1117 => x"536c323a",
  1118 => x"20455345",
  1119 => x"2d52414d",
  1120 => x"20314d42",
  1121 => x"2f415343",
  1122 => x"49493136",
  1123 => x"00000000",
  1124 => x"536c313a",
  1125 => x"204e6f6e",
  1126 => x"65000000",
  1127 => x"536c313a",
  1128 => x"20455345",
  1129 => x"2d534343",
  1130 => x"20314d42",
  1131 => x"2f534343",
  1132 => x"2d490000",
  1133 => x"536c313a",
  1134 => x"204d6567",
  1135 => x"6152414d",
  1136 => x"00000000",
  1137 => x"56474120",
  1138 => x"2d203331",
  1139 => x"4b487a2c",
  1140 => x"20363048",
  1141 => x"7a000000",
  1142 => x"56474120",
  1143 => x"2d203331",
  1144 => x"4b487a2c",
  1145 => x"20353048",
  1146 => x"7a000000",
  1147 => x"5456202d",
  1148 => x"20343830",
  1149 => x"692c2036",
  1150 => x"30487a00",
  1151 => x"496e6974",
  1152 => x"69616c69",
  1153 => x"7a696e67",
  1154 => x"20534420",
  1155 => x"63617264",
  1156 => x"0a000000",
  1157 => x"53444843",
  1158 => x"20636172",
  1159 => x"64206465",
  1160 => x"74656374",
  1161 => x"65640a00",
  1162 => x"46617433",
  1163 => x"32206e6f",
  1164 => x"74207375",
  1165 => x"70706f72",
  1166 => x"7465640a",
  1167 => x"00000000",
  1168 => x"54727969",
  1169 => x"6e672053",
  1170 => x"50454343",
  1171 => x"592e524f",
  1172 => x"4d0a0000",
  1173 => x"53504543",
  1174 => x"43592020",
  1175 => x"524f4d00",
  1176 => x"4c6f6164",
  1177 => x"696e6720",
  1178 => x"42494f53",
  1179 => x"0a000000",
  1180 => x"52656164",
  1181 => x"20666169",
  1182 => x"6c65640a",
  1183 => x"00000000",
  1184 => x"4c6f6164",
  1185 => x"696e6720",
  1186 => x"42494f53",
  1187 => x"20646f6e",
  1188 => x"650a0000",
  1189 => x"4c6f6164",
  1190 => x"696e6720",
  1191 => x"42494f53",
  1192 => x"20666169",
  1193 => x"6c65640a",
  1194 => x"00000000",
  1195 => x"4d425220",
  1196 => x"6661696c",
  1197 => x"0a000000",
  1198 => x"46415431",
  1199 => x"36202020",
  1200 => x"00000000",
  1201 => x"46415433",
  1202 => x"32202020",
  1203 => x"00000000",
  1204 => x"4e6f2070",
  1205 => x"61727469",
  1206 => x"74696f6e",
  1207 => x"20736967",
  1208 => x"0a000000",
  1209 => x"42616420",
  1210 => x"70617274",
  1211 => x"0a000000",
  1212 => x"53444843",
  1213 => x"20657272",
  1214 => x"6f72210a",
  1215 => x"00000000",
  1216 => x"53442069",
  1217 => x"6e69742e",
  1218 => x"2e2e0a00",
  1219 => x"53442063",
  1220 => x"61726420",
  1221 => x"72657365",
  1222 => x"74206661",
  1223 => x"696c6564",
  1224 => x"210a0000",
  1225 => x"57726974",
  1226 => x"65206661",
  1227 => x"696c6564",
  1228 => x"0a000000",
  1229 => x"16200000",
  1230 => x"14200000",
  1231 => x"15200000",
  1232 => x"00000002",
  1233 => x"00000005",
  1234 => x"0000108c",
  1235 => x"00000007",
  1236 => x"00000005",
  1237 => x"00001094",
  1238 => x"00000007",
  1239 => x"00000005",
  1240 => x"0000109c",
  1241 => x"00000007",
  1242 => x"00000005",
  1243 => x"000010a0",
  1244 => x"00000007",
  1245 => x"00000004",
  1246 => x"000010a4",
  1247 => x"0000138c",
  1248 => x"00000000",
  1249 => x"00000000",
  1250 => x"00000000",
  1251 => x"00000002",
  1252 => x"000010ac",
  1253 => x"00000463",
  1254 => x"00000002",
  1255 => x"000010b4",
  1256 => x"00000455",
  1257 => x"00000004",
  1258 => x"000010c4",
  1259 => x"000013ec",
  1260 => x"00000004",
  1261 => x"000010d0",
  1262 => x"00001344",
  1263 => x"00000001",
  1264 => x"000010d8",
  1265 => x"00000007",
  1266 => x"00000001",
  1267 => x"000010e0",
  1268 => x"0000000a",
  1269 => x"00000002",
  1270 => x"000010f0",
  1271 => x"00000f8b",
  1272 => x"00000000",
  1273 => x"00000000",
  1274 => x"00000000",
  1275 => x"00000003",
  1276 => x"0000147c",
  1277 => x"00000003",
  1278 => x"00000001",
  1279 => x"000010f8",
  1280 => x"0000000b",
  1281 => x"00000001",
  1282 => x"00001104",
  1283 => x"00000002",
  1284 => x"00000003",
  1285 => x"00001470",
  1286 => x"00000003",
  1287 => x"00000003",
  1288 => x"00001460",
  1289 => x"00000004",
  1290 => x"00000001",
  1291 => x"0000110c",
  1292 => x"00000006",
  1293 => x"00000003",
  1294 => x"00001458",
  1295 => x"00000002",
  1296 => x"00000004",
  1297 => x"000010a4",
  1298 => x"0000138c",
  1299 => x"00000000",
  1300 => x"00000000",
  1301 => x"00000000",
  1302 => x"00001120",
  1303 => x"0000112c",
  1304 => x"00001138",
  1305 => x"00001144",
  1306 => x"0000115c",
  1307 => x"00001174",
  1308 => x"00001190",
  1309 => x"0000119c",
  1310 => x"000011b4",
  1311 => x"000011c4",
  1312 => x"000011d8",
  1313 => x"000011ec",
  1314 => x"00000003",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

